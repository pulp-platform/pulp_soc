// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.


`include "pulp_soc_defines.sv"
`include "soc_bus_defines.sv"

module pulp_soc import dm::*; #(
    parameter CORE_TYPE          = 0,
    parameter USE_FPU            = 1,
    parameter USE_HWPE           = 1,
    parameter USE_CLUSTER_EVENT  = 1,
    parameter AXI_ADDR_WIDTH     = 32,
    parameter AXI_DATA_IN_WIDTH  = 64,
    parameter AXI_DATA_OUT_WIDTH = 32,
    parameter AXI_ID_IN_WIDTH    = 6,
    parameter AXI_ID_OUT_WIDTH   = 6,
    parameter AXI_USER_WIDTH     = 6,
    parameter AXI_STRB_WIDTH_IN  = AXI_DATA_IN_WIDTH/8,
    parameter AXI_STRB_WIDTH_OUT = AXI_DATA_OUT_WIDTH/8,
    parameter BUFFER_WIDTH       = 8,
    parameter EVNT_WIDTH         = 8,
    parameter NB_CORES           = 8,
    parameter NB_HWPE_PORTS      = 4,
    parameter NGPIO              = 43,
    parameter NPAD               = 64,

    parameter int unsigned AXI_ID_INP_WIDTH_C07 = 6,
    parameter int unsigned AXI_ID_OUP_WIDTH_C07 = 6,
    parameter int unsigned AXI_USER_WIDTH_C07 = 6,
    parameter int unsigned AXI_STRB_WIDTH_C07 = 64/8,
    parameter int unsigned AXI_ADDR_WIDTH_C07 = 32,
    parameter int unsigned AXI_DATA_WIDTH_C07 = 64,

    parameter int unsigned AXI_ID_INP_WIDTH_NOCR07 = 6,
    parameter int unsigned AXI_ID_OUP_WIDTH_NOCR07 = 6,
    parameter int unsigned AXI_USER_WIDTH_NOCR07 = 6,
    parameter int unsigned AXI_STRB_WIDTH_NOCR07 = 64/8,
    parameter int unsigned AXI_ADDR_WIDTH_NOCR07 = 32,
    parameter int unsigned AXI_DATA_WIDTH_NOCR07 = 64,

    parameter int unsigned AXI_ID_WIDTH_SMS = 6,
    parameter int unsigned AXI_USER_WIDTH_SMS = 6,
    parameter int unsigned AXI_STRB_WIDTH_SMS = 64/8,
    parameter int unsigned AXI_ADDR_WIDTH_SMS = 32,
    parameter int unsigned AXI_DATA_WIDTH_SMS = 64,

    parameter NBIT_PADCFG        = 4,
    parameter NBIT_PADMUX        = 2,

    parameter int unsigned N_UART = 1,
    parameter int unsigned N_SPI  = 1,
    parameter int unsigned N_I2C  = 2

) (
    input  logic                          ref_clk_i,
    input  logic                          slow_clk_i,
    input  logic                          test_clk_i,
    input  logic                          rstn_glob_i,

    input  logic                          dft_test_mode_i,
    input  logic                          dft_cg_enable_i,
    input  logic                          mode_select_i,
    input  logic                          boot_l2_i,
    input  logic                          bootsel_i,

    // AXI interfaces to outside of control pulp
    AXI_BUS.Slave                         axi_c07_slv,  // from c07
    AXI_BUS.Master                        axi_c07_mst,

    AXI_BUS.Slave                         axi_nocr07_slv, // from NoC
    AXI_BUS.Master                        axi_nocr07_mst,

    AXI_BUS.Slave                         axi_sms_slv,   // from security subsystem

    output logic                          cluster_rtc_o,
    output logic                          cluster_fetch_enable_o,
    output logic [63:0]                   cluster_boot_addr_o,
    output logic                          cluster_test_en_o,
    output logic                          cluster_pow_o,
    output logic                          cluster_byp_o,
    output logic                          cluster_rstn_o,
    output logic                          cluster_irq_o,
    // AXI4 SLAVE
    input  logic [7:0]                    data_slave_aw_writetoken_i,
    input  logic [AXI_ADDR_WIDTH-1:0]     data_slave_aw_addr_i,
    input  logic [2:0]                    data_slave_aw_prot_i,
    input  logic [3:0]                    data_slave_aw_region_i,
    input  logic [7:0]                    data_slave_aw_len_i,
    input  logic [2:0]                    data_slave_aw_size_i,
    //input  logic [5:0]                    data_slave_aw_atop_i,
    input  logic [1:0]                    data_slave_aw_burst_i,
    input  logic                          data_slave_aw_lock_i,
    input  logic [3:0]                    data_slave_aw_cache_i,
    input  logic [3:0]                    data_slave_aw_qos_i,
    input  logic [AXI_ID_IN_WIDTH-1:0]    data_slave_aw_id_i,
    input  logic [AXI_USER_WIDTH-1:0]     data_slave_aw_user_i,
    output logic [7:0]                    data_slave_aw_readpointer_o,
    input  logic [7:0]                    data_slave_ar_writetoken_i,
    input  logic [AXI_ADDR_WIDTH-1:0]     data_slave_ar_addr_i,
    input  logic [2:0]                    data_slave_ar_prot_i,
    input  logic [3:0]                    data_slave_ar_region_i,
    input  logic [7:0]                    data_slave_ar_len_i,
    input  logic [2:0]                    data_slave_ar_size_i,
    input  logic [1:0]                    data_slave_ar_burst_i,
    input  logic                          data_slave_ar_lock_i,
    input  logic [3:0]                    data_slave_ar_cache_i,
    input  logic [3:0]                    data_slave_ar_qos_i,
    input  logic [AXI_ID_IN_WIDTH-1:0]    data_slave_ar_id_i,
    input  logic [AXI_USER_WIDTH-1:0]     data_slave_ar_user_i,
    output logic [7:0]                    data_slave_ar_readpointer_o,
    input  logic [7:0]                    data_slave_w_writetoken_i,
    input  logic [AXI_DATA_IN_WIDTH-1:0]  data_slave_w_data_i,
    input  logic [AXI_STRB_WIDTH_IN-1:0]  data_slave_w_strb_i,
    input  logic [AXI_USER_WIDTH-1:0]     data_slave_w_user_i,
    input  logic                          data_slave_w_last_i,
    output logic [7:0]                    data_slave_w_readpointer_o,
    output logic [7:0]                    data_slave_r_writetoken_o,
    output logic [AXI_DATA_IN_WIDTH-1:0]  data_slave_r_data_o,
    output logic [1:0]                    data_slave_r_resp_o,
    output logic                          data_slave_r_last_o,
    output logic [AXI_ID_IN_WIDTH-1:0]    data_slave_r_id_o,
    output logic [AXI_USER_WIDTH-1:0]     data_slave_r_user_o,
    input  logic [7:0]                    data_slave_r_readpointer_i,
    output logic [7:0]                    data_slave_b_writetoken_o,
    output logic [1:0]                    data_slave_b_resp_o,
    output logic [AXI_ID_IN_WIDTH-1:0]    data_slave_b_id_o,
    output logic [AXI_USER_WIDTH-1:0]     data_slave_b_user_o,
    input  logic [7:0]                    data_slave_b_readpointer_i,

    // AXI4 MASTER
    output logic [7:0]                    data_master_aw_writetoken_o,
    output logic [AXI_ADDR_WIDTH-1:0]     data_master_aw_addr_o,
    output logic [2:0]                    data_master_aw_prot_o,
    output logic [3:0]                    data_master_aw_region_o,
    output logic [7:0]                    data_master_aw_len_o,
    output logic [2:0]                    data_master_aw_size_o,
    // output logic [5:0]                    data_master_aw_atop_o,
    output logic [1:0]                    data_master_aw_burst_o,
    output logic                          data_master_aw_lock_o,
    output logic [3:0]                    data_master_aw_cache_o,
    output logic [3:0]                    data_master_aw_qos_o,
    output logic [AXI_ID_OUT_WIDTH-1:0]   data_master_aw_id_o,
    output logic [AXI_USER_WIDTH-1:0]     data_master_aw_user_o,
    input  logic [7:0]                    data_master_aw_readpointer_i,
    output logic [7:0]                    data_master_ar_writetoken_o,
    output logic [AXI_ADDR_WIDTH-1:0]     data_master_ar_addr_o,
    output logic [2:0]                    data_master_ar_prot_o,
    output logic [3:0]                    data_master_ar_region_o,
    output logic [7:0]                    data_master_ar_len_o,
    output logic [2:0]                    data_master_ar_size_o,
    output logic [1:0]                    data_master_ar_burst_o,
    output logic                          data_master_ar_lock_o,
    output logic [3:0]                    data_master_ar_cache_o,
    output logic [3:0]                    data_master_ar_qos_o,
    output logic [AXI_ID_OUT_WIDTH-1:0]   data_master_ar_id_o,
    output logic [AXI_USER_WIDTH-1:0]     data_master_ar_user_o,
    input  logic [7:0]                    data_master_ar_readpointer_i,
    output logic [7:0]                    data_master_w_writetoken_o,
    output logic [AXI_DATA_OUT_WIDTH-1:0] data_master_w_data_o,
    output logic [AXI_STRB_WIDTH_OUT-1:0] data_master_w_strb_o,
    output logic [AXI_USER_WIDTH-1:0]     data_master_w_user_o,
    output logic                          data_master_w_last_o,
    input  logic [7:0]                    data_master_w_readpointer_i,
    input  logic [7:0]                    data_master_r_writetoken_i,
    input  logic [AXI_DATA_OUT_WIDTH-1:0] data_master_r_data_i,
    input  logic [1:0]                    data_master_r_resp_i,
    input  logic                          data_master_r_last_i,
    input  logic [AXI_ID_OUT_WIDTH-1:0]   data_master_r_id_i,
    input  logic [AXI_USER_WIDTH-1:0]     data_master_r_user_i,
    output logic [7:0]                    data_master_r_readpointer_o,
    input  logic [7:0]                    data_master_b_writetoken_i,
    input  logic [1:0]                    data_master_b_resp_i,
    input  logic [AXI_ID_OUT_WIDTH-1:0]   data_master_b_id_i,
    input  logic [AXI_USER_WIDTH-1:0]     data_master_b_user_i,
    output logic [7:0]                    data_master_b_readpointer_o,

    output logic [BUFFER_WIDTH-1:0]       cluster_events_wt_o,
    input  logic [BUFFER_WIDTH-1:0]       cluster_events_rp_i,
    output logic [EVNT_WIDTH-1:0]         cluster_events_da_o,
    output logic                          cluster_clk_o,
    input  logic                          cluster_busy_i,
    output logic                          dma_pe_evt_ack_o,
    input  logic                          dma_pe_evt_valid_i,
    output logic                          dma_pe_irq_ack_o,
    input  logic                          dma_pe_irq_valid_i,
    output logic                          pf_evt_ack_o,
    input  logic                          pf_evt_valid_i,
    ///////////////////////////////////////////////////
    //      To I/O Controller and padframe           //
    ///////////////////////////////////////////////////
    output logic [127:0]                  pad_mux_o,
    output logic [383:0]                  pad_cfg_o,
    input  logic [31:0]                   gpio_in_i,
    output logic [31:0]                   gpio_out_o,
    output logic [31:0]                   gpio_dir_o,
    output logic [191:0]                  gpio_cfg_o,
    output logic                          uart_tx_o,
    input  logic                          uart_rx_i,
    input  logic                          cam_clk_i,
    input  logic [7:0]                    cam_data_i,
    input  logic                          cam_hsync_i,
    input  logic                          cam_vsync_i,
    output logic [3:0]                    timer_ch0_o,
    output logic [3:0]                    timer_ch1_o,
    output logic [3:0]                    timer_ch2_o,
    output logic [3:0]                    timer_ch3_o,

    // input  logic                          i2c0_scl_i,
    // output logic                          i2c0_scl_o,
    // output logic                          i2c0_scl_oe_o,
    // input  logic                          i2c0_sda_i,
    // output logic                          i2c0_sda_o,
    // output logic                          i2c0_sda_oe_o,
    // input  logic                          i2c1_scl_i,
    // output logic                          i2c1_scl_o,
    // output logic                          i2c1_scl_oe_o,
    // input  logic                          i2c1_sda_i,
    // output logic                          i2c1_sda_o,
    // output logic                          i2c1_sda_oe_o,

    input  logic [N_I2C-1:0]              i2c_scl_i,
    output logic [N_I2C-1:0]              i2c_scl_o,
    output logic [N_I2C-1:0]              i2c_scl_oe_o,
    input  logic [N_I2C-1:0]              i2c_sda_i,
    output logic [N_I2C-1:0]              i2c_sda_o,
    output logic [N_I2C-1:0]              i2c_sda_oe_o,

    input  logic                          i2s_slave_sd0_i,
    input  logic                          i2s_slave_sd1_i,
    input  logic                          i2s_slave_ws_i,
    output logic                          i2s_slave_ws_o,
    output logic                          i2s_slave_ws_oe,
    input  logic                          i2s_slave_sck_i,
    output logic                          i2s_slave_sck_o,
    output logic                          i2s_slave_sck_oe,
    output logic                          spi_master0_clk_o,
    output logic                          spi_master0_csn0_o,
    output logic                          spi_master0_csn1_o,
    output logic                          spi_master0_oen0_o,
    output logic                          spi_master0_oen1_o,
    output logic                          spi_master0_oen2_o,
    output logic                          spi_master0_oen3_o,
    output logic                          spi_master0_sdo0_o,
    output logic                          spi_master0_sdo1_o,
    output logic                          spi_master0_sdo2_o,
    output logic                          spi_master0_sdo3_o,
    input  logic                          spi_master0_sdi0_i,
    input  logic                          spi_master0_sdi1_i,
    input  logic                          spi_master0_sdi2_i,
    input  logic                          spi_master0_sdi3_i,
    output logic                          sdio_clk_o,
    output logic                          sdio_cmd_o,
    input  logic                          sdio_cmd_i,
    output logic                          sdio_cmd_oen_o,
    output logic                    [3:0] sdio_data_o,
    input  logic                    [3:0] sdio_data_i,
    output logic                    [3:0] sdio_data_oen_o,

    ///////////////////////////////////////////////////
    ///////////////////////////////////////////////////
    // From JTAG Tap Controller to axi_dcb module    //
    ///////////////////////////////////////////////////
    input  logic                          jtag_tck_i,
    input  logic                          jtag_trst_ni,
    input  logic                          jtag_tms_i,
    input  logic                          jtag_tdi_i,
    output logic                          jtag_tdo_o,
    output logic [NB_CORES-1:0]          cluster_dbg_irq_valid_o
    ///////////////////////////////////////////////////
);

    genvar dbg_var, nhart_var;

    localparam FLL_ADDR_WIDTH        = 32;
    localparam FLL_DATA_WIDTH        = 32;
    localparam NB_L2_BANKS           = `NB_L2_CHANNELS;
    localparam L2_BANK_SIZE          = 29184;            // in 32-bit words
    localparam L2_MEM_ADDR_WIDTH     = $clog2(L2_BANK_SIZE * NB_L2_BANKS) - $clog2(NB_L2_BANKS);    // 2**L2_MEM_ADDR_WIDTH rows (64bit each) in L2 --> TOTAL L2 SIZE = 8byte * 2^L2_MEM_ADDR_WIDTH
    localparam NB_L2_BANKS_PRI       = 2;
    localparam L2_BANK_SIZE_PRI      = 8192;             // in 32-bit words
    localparam L2_MEM_ADDR_WIDTH_PRI = $clog2(L2_BANK_SIZE_PRI * NB_L2_BANKS_PRI) - $clog2(NB_L2_BANKS_PRI);
    localparam ROM_ADDR_WIDTH        = 13;

    localparam FC_Core_CLUSTER_ID    = 6'd31;
    localparam CL_Core_CLUSTER_ID    = 6'd0;

    localparam FC_Core_CORE_ID       = 4'd0;
    localparam FC_Core_MHARTID       = {FC_Core_CLUSTER_ID,1'b0,FC_Core_CORE_ID};
    localparam CL_Core0_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd0};
    localparam CL_Core1_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd1};
    localparam CL_Core2_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd2};
    localparam CL_Core3_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd3};
    localparam CL_Core4_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd4};
    localparam CL_Core5_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd5};
    localparam CL_Core6_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd6};
    localparam CL_Core7_MHARTID      = {CL_Core_CLUSTER_ID,1'b0,4'd7};


    // TODO: this should be exposed somewhere, maybe configurable?
    localparam int unsigned AXI_SOC_NODE_AW = 32;
    localparam int unsigned AXI_SOC_NODE_DW = 64;
    localparam int unsigned AXI_SOC_NODE_UW = 6;
    localparam int unsigned AXI_SOC_NODE_IW_INP = 6;
    localparam int unsigned AXI_SOC_NODE_IW_OUP = soc_node_pkg::axi_iw_oup(AXI_SOC_NODE_IW_INP);

    /*
        PULP RISC-V cores have not continguos MHARTID.
        This leads to set the number of HARTS >= the maximum value of the MHARTID.
        In this case, the MHARD ID is {FC_Core_CLUSTER_ID,1'b0,FC_Core_CORE_ID} --> 996 (1024 chosen as power of 2)
        To avoid paying 1024 flip flop for each number of harts's related register, we implemented
        the masking parameter, aka SELECTABLE_HARTS.
        In One-Hot-Encoding way, you select 1 when that MHARTID-related HART can actally be selected.
        e.g. if you have 2 core with MHART 10 and 5, you select NrHarts=16 and SELECTABLE_HARTS = (1<<10) | (1<<5).
        This mask will be used to generated only the flip flop needed and the constant-propagator engine of the synthesizer
        will remove the other flip flops and related logic.
    */

    localparam NrHarts                               = 1024;
    localparam logic [NrHarts-1:0] SELECTABLE_HARTS  = (1 << FC_Core_MHARTID) | (1 << CL_Core0_MHARTID) | (1 << CL_Core1_MHARTID) | (1 << CL_Core2_MHARTID) | (1 << CL_Core3_MHARTID) | (1 << CL_Core4_MHARTID) | (1 << CL_Core5_MHARTID) | (1 << CL_Core6_MHARTID) | (1 << CL_Core7_MHARTID);

    logic [NB_CORES-1:0][10:0]   CLUSTER_CORE_ID;

    assign CLUSTER_CORE_ID[0] = CL_Core0_MHARTID;
    assign CLUSTER_CORE_ID[1] = CL_Core1_MHARTID;
    assign CLUSTER_CORE_ID[2] = CL_Core2_MHARTID;
    assign CLUSTER_CORE_ID[3] = CL_Core3_MHARTID;
    assign CLUSTER_CORE_ID[4] = CL_Core4_MHARTID;
    assign CLUSTER_CORE_ID[5] = CL_Core5_MHARTID;
    assign CLUSTER_CORE_ID[6] = CL_Core6_MHARTID;
    assign CLUSTER_CORE_ID[7] = CL_Core7_MHARTID;


    localparam dm::hartinfo_t RI5CY_HARTINFO = '{
                                                zero1:        '0,
                                                nscratch:      2, // Debug module needs at least two scratch regs
                                                zero0:        '0,
                                                dataaccess: 1'b1, // data registers are memory mapped in the debugger
                                                datasize: dm::DataCount,
                                                dataaddr: dm::DataAddr
                                               };

    dm::hartinfo_t [NrHarts-1:0] hartinfo;

    /*
       This module has been tested only with the default parameters.
    */

    //********************************************************
    //***************** SIGNALS DECLARATION ******************
    //********************************************************
    logic [ 1:0]           s_fc_hwpe_events;
    logic [31:0]           s_fc_events;

    logic [7:0]            s_soc_events_ack;
    logic [7:0]            s_soc_events_val;

    logic                  s_timer_lo_event;
    logic                  s_timer_hi_event;

    logic [EVNT_WIDTH-1:0] s_cl_event_data ;
    logic                  s_cl_event_valid;
    logic                  s_cl_event_ready;

    logic [EVNT_WIDTH-1:0] s_fc_event_data ;
    logic                  s_fc_event_valid;
    logic                  s_fc_event_ready;

    logic [7:0][31:0]      s_apb_mpu_rules;
    logic                  s_supervisor_mode;

    logic [31:0]           s_fc_bootaddr;

    logic [31:0][5:0]      s_gpio_cfg;
    logic [63:0][1:0]      s_pad_mux;
    logic [63:0][5:0]      s_pad_cfg;

    logic                  s_periph_clk;
    logic                  s_periph_rstn;
    logic                  s_soc_clk;
    logic                  s_soc_rstn;
    logic                  s_cluster_clk;
    logic                  s_cluster_rstn;
    logic                  s_cluster_rstn_soc_ctrl;
    logic                  s_sel_fll_clk;

    logic                  s_dma_pe_evt;
    logic                  s_dma_pe_irq;
    logic                  s_pf_evt;

    logic                  s_fc_fetchen;
    logic [NrHarts-1:0]    dm_debug_req;

    logic                  jtag_req_valid;
    logic                  debug_req_ready;
    logic                  jtag_resp_ready;
    logic                  jtag_resp_valid;
    dm::dmi_req_t          jtag_dmi_req;
    dm::dmi_resp_t         debug_resp;
    logic                  slave_grant, slave_valid, slave_req , slave_we;
    logic                  [31:0] slave_addr, slave_wdata, slave_rdata;
    logic                  [3:0]  slave_be;
    logic                  lint_riscv_jtag_bus_master_we;
    logic                  int_td;

    logic                  master_req;
    logic [31:0]           master_add;
    logic                  master_we;
    logic [31:0]           master_wdata;
    logic [3:0]            master_be;
    logic                  master_gnt;
    logic                  master_r_valid;
    logic [31:0]           master_r_rdata;


    logic [7:0]            soc_jtag_reg_tap;
    logic [7:0]            soc_jtag_reg_soc;


    logic                  spi_master0_csn3, spi_master0_csn2;

    genvar                 i,j;

    //wdt reset output:
    logic			wdt_reset_o;

    APB_BUS                s_apb_eu_bus ();
    APB_BUS                s_apb_hwpe_bus ();
    APB_BUS                s_apb_debug_bus();

    AXI_BUS_ASYNC #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_OUT_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     ),
        .BUFFER_WIDTH   ( BUFFER_WIDTH       )
    ) s_data_master ();

    AXI_BUS_ASYNC #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    ),
        .BUFFER_WIDTH   ( BUFFER_WIDTH      )
    ) s_data_slave ();

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_data_in_bus ();

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_WIDTH),
        .AXI_ID_WIDTH   ( AXI_ID_OUT_WIDTH  ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_data_out_bus ();

    // cl master -> soc_node
    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_OUT_WIDTH  ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) cl_in_mst ();

    // soc_node -> soc
    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH      ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH   ),
        .AXI_ID_WIDTH   ( AXI_SOC_NODE_IW_OUP ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH      )
    ) soc_in_mst ();

    //assign s_data_out_bus.aw_atop = 6'b0;

    FLL_BUS #(
        .FLL_ADDR_WIDTH ( FLL_ADDR_WIDTH ),
        .FLL_DATA_WIDTH ( FLL_DATA_WIDTH )
    ) s_soc_fll_master ();

    FLL_BUS #(
        .FLL_ADDR_WIDTH ( FLL_ADDR_WIDTH ),
        .FLL_DATA_WIDTH ( FLL_DATA_WIDTH )
    ) s_per_fll_master ();

    FLL_BUS #(
        .FLL_ADDR_WIDTH ( FLL_ADDR_WIDTH ),
        .FLL_DATA_WIDTH ( FLL_DATA_WIDTH )
    ) s_cluster_fll_master ();

    APB_BUS s_apb_periph_bus ();

    UNICAD_MEM_BUS_32 s_mem_rom_bus ();

    UNICAD_MEM_BUS_32  s_mem_l2_bus[NB_L2_BANKS-1:0]();
    UNICAD_MEM_BUS_32  s_mem_l2_pri_bus[NB_L2_BANKS_PRI-1:0]();
`ifdef QUENTIN_SCM
    UNICAD_MEM_BUS_32 s_scm_l2_data_bus ();
    UNICAD_MEM_BUS_32 s_scm_l2_instr_bus ();
`endif

    XBAR_TCDM_BUS s_lint_debug_bus();
    XBAR_TCDM_BUS s_lint_pulp_jtag_bus();
    XBAR_TCDM_BUS s_lint_riscv_jtag_bus();
    XBAR_TCDM_BUS s_lint_udma_tx_bus ();
    XBAR_TCDM_BUS s_lint_udma_rx_bus ();
    XBAR_TCDM_BUS s_lint_fc_data_bus ();
    XBAR_TCDM_BUS s_lint_fc_instr_bus ();
    XBAR_TCDM_BUS s_lint_hwpe_bus[NB_HWPE_PORTS-1:0]();

    `ifdef REMAP_ADDRESS
        logic [3:0] base_addr_int;
        assign base_addr_int = 4'b0001; //FIXME attach this signal somewhere in the soc peripherals --> IGOR
    `endif



    logic s_cluster_isolate_dc;
    logic s_rstn_cluster_sync_soc;


    assign cluster_clk_o  = s_cluster_clk;
    assign cluster_rstn_o = s_cluster_rstn && s_cluster_rstn_soc_ctrl;
    assign s_rstn_cluster_sync_soc = s_cluster_rstn && s_cluster_rstn_soc_ctrl;

    assign cluster_rtc_o     = ref_clk_i;
    assign cluster_test_en_o = dft_test_mode_i;
    // isolate dc if the cluster is down
   assign s_cluster_isolate_dc = 1'b0;
//cluster_byp_o;
    // If you want to connect a real PULP cluster you also need a cluster_busy_i signal

    // cluster to soc
    axi_slice_dc_master_wrap  #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    ),
        .BUFFER_WIDTH   ( BUFFER_WIDTH      )
    ) dc_fifo_dataout_bus_i (
        .clk_i           ( s_soc_clk                ),
        .rst_ni          ( s_cluster_rstn           ),
        .isolate_i       ( s_cluster_isolate_dc     ),
        .test_cgbypass_i ( 1'b0                     ),
        .clock_down_i    ( 1'b0                     ),
        .incoming_req_o  (                          ),
        .axi_master      ( s_data_in_bus            ),
        .axi_slave_async ( s_data_slave             )
    );

    // soc to cluster
    axi_slice_dc_slave_wrap #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_OUT_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     ),
        .BUFFER_WIDTH   ( BUFFER_WIDTH       )
    ) dc_fifo_datain_bus_i (
        .clk_i            ( s_soc_clk               ),
        .rst_ni           ( s_rstn_cluster_sync_soc ),
        .test_cgbypass_i  ( 1'b0                    ),
        .isolate_i        ( s_cluster_isolate_dc    ),
        .axi_slave        ( s_data_out_bus          ),
        .axi_master_async ( s_data_master           )
    );


    // data width conversions of AXI to 32-bit. Currently we fail here if we have
    // a mismatch.
    if (AXI_DATA_IN_WIDTH != AXI_DATA_WIDTH_C07)
        $fatal("AXI data width mismatch on c07");
    if (AXI_DATA_IN_WIDTH != AXI_DATA_WIDTH_NOCR07)
        $fatal("AXI data width mismatch on nocr07");
    if (AXI_DATA_IN_WIDTH != AXI_DATA_WIDTH_SMS)
        $fatal("AXI data width mismatch on sms");
    /* axi_data_width_converter AUTO_TEMPLATE "_\([a-z]+\)" (
     .slv (axi_in[]),
     .mst (axi[]),
     );
     */

    // Addr width conversion of AXI. Currently we fail here if we have a mismatch.
    if (AXI_ADDR_WIDTH != AXI_ADDR_WIDTH_C07)
        $fatal("AXI address width mismatch on c07");
    if (AXI_ADDR_WIDTH != AXI_ADDR_WIDTH_NOCR07)
        $fatal("AXI address width mismatch on nocr07");
    if (AXI_ADDR_WIDTH != AXI_ADDR_WIDTH_SMS)
        $fatal("AXI address width mismatch on sms");

    //
    // AXI soc node
    //
    // We connect the axi bus from the cluster with all the external axi master
    // and slaves and route this to the tcdm interconnect

    soc_node #(
        // Parameters
        .AXI_ID_OUP_WIDTH_SOC    (AXI_SOC_NODE_IW_OUP),
        .AXI_USER_WIDTH_SOC      (AXI_USER_WIDTH),
        .AXI_STRB_WIDTH_SOC      (AXI_DATA_IN_WIDTH/8),
        .AXI_ADDR_WIDTH_SOC      (AXI_ADDR_WIDTH),
        .AXI_DATA_WIDTH_SOC      (AXI_DATA_IN_WIDTH),

        .AXI_ID_INP_WIDTH_CLUSTER(AXI_ID_IN_WIDTH),
        .AXI_USER_WIDTH_CLUSTER  (AXI_USER_WIDTH),
        .AXI_STRB_WIDTH_CLUSTER  (AXI_DATA_IN_WIDTH/8),
        .AXI_ADDR_WIDTH_CLUSTER  (AXI_ADDR_WIDTH),
        .AXI_DATA_WIDTH_CLUSTER  (AXI_DATA_IN_WIDTH),

        .AXI_ID_INP_WIDTH_C07    (AXI_ID_INP_WIDTH_C07),
        .AXI_ID_OUP_WIDTH_C07    (AXI_ID_OUP_WIDTH_C07),
        .AXI_USER_WIDTH_C07      (AXI_USER_WIDTH_C07),
        .AXI_STRB_WIDTH_C07      (AXI_STRB_WIDTH_C07),
        .AXI_ADDR_WIDTH_C07      (AXI_ADDR_WIDTH_C07),
        .AXI_DATA_WIDTH_C07      (AXI_DATA_WIDTH_C07),

        .AXI_ID_INP_WIDTH_NOCR07 (AXI_ID_INP_WIDTH_NOCR07),
        .AXI_ID_OUP_WIDTH_NOCR07 (AXI_ID_OUP_WIDTH_NOCR07),
        .AXI_USER_WIDTH_NOCR07   (AXI_USER_WIDTH_NOCR07),
        .AXI_STRB_WIDTH_NOCR07   (AXI_STRB_WIDTH_NOCR07),
        .AXI_ADDR_WIDTH_NOCR07   (AXI_ADDR_WIDTH_NOCR07),
        .AXI_DATA_WIDTH_NOCR07   (AXI_DATA_WIDTH_NOCR07),

        .AXI_ID_INP_WIDTH_SMS    (AXI_ID_WIDTH_SMS),
        .AXI_USER_WIDTH_SMS      (AXI_USER_WIDTH_SMS),
        .AXI_STRB_WIDTH_SMS      (AXI_STRB_WIDTH_SMS),
        .AXI_ADDR_WIDTH_SMS      (AXI_ADDR_WIDTH_SMS),
        .AXI_DATA_WIDTH_SMS      (AXI_DATA_WIDTH_SMS),

        // this is the soc nodes axi config. All connections' parameters will be
        // checked against this
        .AXI_AW                  (AXI_SOC_NODE_AW),
        .AXI_DW                  (AXI_SOC_NODE_DW),
        .AXI_UW                  (AXI_SOC_NODE_UW),
        .AXI_IW_INP              (AXI_SOC_NODE_IW_INP), // cluster -> soc id width
        .MST_SLICE_DEPTH         (1),
        .SLV_SLICE_DEPTH         (1)
    ) i_soc_node (
        // Interfaces
        .cl_slv          (s_data_in_bus),
        //.cl_mst          (cl_in_Mst),
        .soc_mst         (soc_in_mst),
        .c07_slv         (axi_c07_slv),
        .c07_mst         (axi_c07_mst),
        .nocr07_slv      (axi_nocr07_slv),
        .nocr07_mst      (axi_nocr07_mst),
        .sms_slv         (axi_sms_slv),
        // Inputs
        .clk_i           (s_soc_clk),
        .rst_ni          (s_soc_rstn)
    );


    //********************************************************
    //********************* SOC L2 RAM ***********************
    //********************************************************

    l2_ram_multi_bank #(
        .MEM_ADDR_WIDTH        ( L2_MEM_ADDR_WIDTH     ),
        .NB_BANKS              ( NB_L2_BANKS           ),
        .BANK_SIZE             ( L2_BANK_SIZE          ),
        .MEM_ADDR_WIDTH_PRI    ( L2_MEM_ADDR_WIDTH_PRI ),
        .NB_BANKS_PRI          ( NB_L2_BANKS_PRI       )
    ) l2_ram_i (
        .clk_i           ( s_soc_clk          ),
        .rst_ni          ( s_soc_rstn         ),
        .init_ni         ( 1'b1               ),
        .test_mode_i     ( dft_test_mode_i    ),
        .mem_slave       ( s_mem_l2_bus       ),
        .mem_pri_slave   ( s_mem_l2_pri_bus   )
`ifdef QUENTIN_SCM
        ,
        .scm_data_slave  ( s_scm_l2_data_bus  ),
        .scm_instr_slave ( s_scm_l2_instr_bus )
`endif
    );


    //********************************************************
    //******              SOC BOOT ROM             ***********
    //********************************************************

    boot_rom #(
        .ROM_ADDR_WIDTH(ROM_ADDR_WIDTH)
    ) boot_rom_i (
        .clk_i       ( s_soc_clk       ),
        .rst_ni      ( s_soc_rstn      ),
        .init_ni     ( 1'b1            ),
        .mem_slave   ( s_mem_rom_bus   ),
        .test_mode_i ( dft_test_mode_i )
    );

    //********************************************************
    //********************* SOC PERIPHERALS ******************
    //********************************************************

    soc_peripherals #(
        .CORE_TYPE          ( CORE_TYPE                             ),
        .MEM_ADDR_WIDTH     ( L2_MEM_ADDR_WIDTH+$clog2(NB_L2_BANKS) ),
        .APB_ADDR_WIDTH     ( 32                                    ),
        .APB_DATA_WIDTH     ( 32                                    ),
        .NB_CORES           ( NB_CORES                              ),
        .NB_CLUSTERS        ( `NB_CLUSTERS                          ),
        .EVNT_WIDTH         ( EVNT_WIDTH                            ),
        .NGPIO              ( NGPIO                                 ),
        .NPAD               ( NPAD                                  ),
        .NBIT_PADCFG        ( NBIT_PADCFG                           ),
        .NBIT_PADMUX        ( NBIT_PADMUX                           ),
        .N_UART             ( N_UART                                ),
        .N_SPI              ( N_SPI                                 ),
        .N_I2C              ( N_I2C                                 )
    ) soc_peripherals_i (

        .clk_i                  ( s_soc_clk              ),
        .periph_clk_i           ( s_periph_clk           ),
        .rst_ni                 ( s_soc_rstn             ),
        .sel_fll_clk_i          ( s_sel_fll_clk          ),
        .ref_clk_i              ( ref_clk_i              ),
        .slow_clk_i             ( slow_clk_i             ),

        .dft_test_mode_i        ( dft_test_mode_i        ),
        .dft_cg_enable_i        ( 1'b0                   ),

        .boot_l2_i              ( boot_l2_i              ),
        .bootsel_i              ( bootsel_i              ),

        .fc_bootaddr_o          ( s_fc_bootaddr          ),
        .fc_fetchen_o           ( s_fc_fetchen           ),

        .apb_slave              ( s_apb_periph_bus       ),

        .apb_eu_master          ( s_apb_eu_bus           ),
        .apb_debug_master       ( s_apb_debug_bus        ),
        .apb_hwpe_master        ( s_apb_hwpe_bus         ),

        .l2_rx_master           ( s_lint_udma_rx_bus     ),
        .l2_tx_master           ( s_lint_udma_tx_bus     ),

        .soc_jtag_reg_i         ( soc_jtag_reg_tap       ),
        .soc_jtag_reg_o         ( soc_jtag_reg_soc       ),

        .fc_hwpe_events_i       ( s_fc_hwpe_events       ),
        .fc_events_o            ( s_fc_events            ),

        .dma_pe_evt_i           ( s_dma_pe_evt           ),
        .dma_pe_irq_i           ( s_dma_pe_irq           ),
        .pf_evt_i               ( s_pf_evt               ),

        .soc_fll_master         ( s_soc_fll_master       ),
        .per_fll_master         ( s_per_fll_master       ),
        .cluster_fll_master     ( s_cluster_fll_master   ),

        .gpio_in                ( gpio_in_i              ),
        .gpio_out               ( gpio_out_o             ),
        .gpio_dir               ( gpio_dir_o             ),
        .gpio_padcfg            ( s_gpio_cfg             ),

        .pad_mux_o              ( s_pad_mux              ),
        .pad_cfg_o              ( s_pad_cfg              ),

        //CAMERA
        .cam_clk_i              ( cam_clk_i              ),
        .cam_data_i             ( cam_data_i             ),
        .cam_hsync_i            ( cam_hsync_i            ),
        .cam_vsync_i            ( cam_vsync_i            ),

        //UART
        .uart_tx                ( uart_tx_o              ),
        .uart_rx                ( uart_rx_i              ),

        //I2C
        .i2c_scl_i              ( i2c_scl_i              ),
        .i2c_scl_o              ( i2c_scl_o              ),
        .i2c_scl_oe_o           ( i2c_scl_oe_o           ),
        .i2c_sda_i              ( i2c_sda_i              ),
        .i2c_sda_o              ( i2c_sda_o              ),
        .i2c_sda_oe_o           ( i2c_sda_oe_o           ),

        //I2S
        .i2s_slave_sd0_i        ( i2s_slave_sd0_i        ),
        .i2s_slave_sd1_i        ( i2s_slave_sd1_i        ),
        .i2s_slave_ws_i         ( i2s_slave_ws_i         ),
        .i2s_slave_ws_o         ( i2s_slave_ws_o         ),
        .i2s_slave_ws_oe        ( i2s_slave_ws_oe        ),
        .i2s_slave_sck_i        ( i2s_slave_sck_i        ),
        .i2s_slave_sck_o        ( i2s_slave_sck_o        ),
        .i2s_slave_sck_oe       ( i2s_slave_sck_oe       ),

         //SPI
        .spi_clk     ( spi_master0_clk_o      ),
        .spi_csn     ( {spi_master0_csn3, spi_master0_csn2, spi_master0_csn1_o, spi_master0_csn0_o}     ), //csn3 and csn2 unconnected
        .spi_oen     ( {spi_master0_oen3_o, spi_master0_oen2_o, spi_master0_oen1_o, spi_master0_oen0_o} ),
        .spi_sdo     ( {spi_master0_sdo3_o, spi_master0_sdo2_o, spi_master0_sdo1_o, spi_master0_sdo0_o} ),
        .spi_sdi     ( {spi_master0_sdi3_i, spi_master0_sdi2_i, spi_master0_sdi1_i, spi_master0_sdi0_i} ),

        //SDIO
        .sdclk_o                ( sdio_clk_o             ),
        .sdcmd_o                ( sdio_cmd_o             ),
        .sdcmd_i                ( sdio_cmd_i             ),
        .sdcmd_oen_o            ( sdio_cmd_oen_o         ),
        .sddata_o               ( sdio_data_o            ),
        .sddata_i               ( sdio_data_i            ),
        .sddata_oen_o           ( sdio_data_oen_o        ),

        .timer_ch0_o            ( timer_ch0_o            ),
        .timer_ch1_o            ( timer_ch1_o            ),
        .timer_ch2_o            ( timer_ch2_o            ),
        .timer_ch3_o            ( timer_ch3_o            ),

        .cl_event_data_o        ( s_cl_event_data        ),
        .cl_event_valid_o       ( s_cl_event_valid       ),
        .cl_event_ready_i       ( s_cl_event_ready       ),

        .fc_event_data_o        ( s_fc_event_data        ),
        .fc_event_valid_o       ( s_fc_event_valid       ),
        .fc_event_ready_i       ( s_fc_event_ready       ),

        .cluster_pow_o          ( cluster_pow_o          ),
        .cluster_byp_o          ( cluster_byp_o          ),
        .cluster_boot_addr_o    ( cluster_boot_addr_o    ),
        .cluster_fetch_enable_o ( cluster_fetch_enable_o ),
        .cluster_rstn_o         ( s_cluster_rstn_soc_ctrl),
        .cluster_irq_o          ( cluster_irq_o          ),

        .wdt_reset_o		( wdt_reset_o		 )
    );



    dc_token_ring_fifo_din #(
        .DATA_WIDTH   ( EVNT_WIDTH   ),
        .BUFFER_DEPTH ( BUFFER_WIDTH )
    ) u_event_dc (
        .clk          ( s_soc_clk               ),
        .rstn         ( s_rstn_cluster_sync_soc ),
        .data         ( s_cl_event_data         ),
        .valid        ( s_cl_event_valid        ),
        .ready        ( s_cl_event_ready        ),
        .write_token  ( cluster_events_wt_o     ),
        .read_pointer ( cluster_events_rp_i     ),
        .data_async   ( cluster_events_da_o     )
    );


    edge_propagator_rx ep_dma_pe_evt_i (
        .clk_i   ( s_soc_clk               ),
        .rstn_i  ( s_rstn_cluster_sync_soc ),
        .valid_o ( s_dma_pe_evt            ),
        .ack_o   ( dma_pe_evt_ack_o        ),
        .valid_i ( dma_pe_evt_valid_i      )
    );

    edge_propagator_rx ep_dma_pe_irq_i (
        .clk_i   ( s_soc_clk               ),
        .rstn_i  ( s_rstn_cluster_sync_soc ),
        .valid_o ( s_dma_pe_irq            ),
        .ack_o   ( dma_pe_irq_ack_o        ),
        .valid_i ( dma_pe_irq_valid_i      )
    );
`ifndef PULP_FPGA_EMUL
    edge_propagator_rx ep_pf_evt_i (
        .clk_i   ( s_soc_clk               ),
        .rstn_i  ( s_rstn_cluster_sync_soc ),
        .valid_o ( s_pf_evt                ),
        .ack_o   ( pf_evt_ack_o            ),
        .valid_i ( pf_evt_valid_i          )
    );
`endif

    fc_subsystem #(
        .CORE_TYPE  ( CORE_TYPE          ),
        .USE_FPU    ( USE_FPU            ),
        .CORE_ID    ( FC_Core_CORE_ID    ),
        .CLUSTER_ID ( FC_Core_CLUSTER_ID ),
        .USE_HWPE   ( USE_HWPE           )
    ) fc_subsystem_i (
        .clk_i               ( s_soc_clk           ),
        .rst_ni              ( s_soc_rstn          ),

        .test_en_i           ( dft_test_mode_i     ),

        //wdt
        .wdt_reset_i	     ( wdt_reset_o         ),

        .boot_addr_i         ( s_fc_bootaddr       ),

        .fetch_en_i          ( s_fc_fetchen        ),

        .l2_data_master      ( s_lint_fc_data_bus  ),
        .l2_instr_master     ( s_lint_fc_instr_bus ),
        .l2_hwpe_master      ( s_lint_hwpe_bus     ),
`ifdef QUENTIN_SCM
        .scm_l2_data_master  ( s_scm_l2_data_bus   ),
        .scm_l2_instr_master ( s_scm_l2_instr_bus  ),
`endif
        .apb_slave_eu        ( s_apb_eu_bus        ),
        .apb_slave_hwpe      ( s_apb_hwpe_bus      ),
        .debug_req_i         ( dm_debug_req[FC_Core_MHARTID] ),

        .event_fifo_valid_i  ( s_fc_event_valid    ),
        .event_fifo_fulln_o  ( s_fc_event_ready    ),
        .event_fifo_data_i   ( s_fc_event_data     ),
        .events_i            ( s_fc_events         ),
        .hwpe_events_o       ( s_fc_hwpe_events    ),

        .supervisor_mode_o   ( s_supervisor_mode   )
    );

    soc_clk_rst_gen i_clk_rst_gen (
        .ref_clk_i                  ( ref_clk_i                     ),
        .test_clk_i                 ( test_clk_i                    ),
        .sel_fll_clk_i              ( s_sel_fll_clk                 ),

        .rstn_glob_i                ( rstn_glob_i                   ),
        .rstn_soc_sync_o            ( s_soc_rstn                    ),
        .rstn_cluster_sync_o        ( s_cluster_rstn                ),

        .clk_cluster_o              ( s_cluster_clk                 ),
        .test_mode_i                ( dft_test_mode_i               ),
        .shift_enable_i             ( 1'b0                          ),

        .soc_fll_slave_req_i        ( s_soc_fll_master.req          ),
        .soc_fll_slave_wrn_i        ( s_soc_fll_master.wrn          ),
        .soc_fll_slave_add_i        ( s_soc_fll_master.add[1:0]     ),
        .soc_fll_slave_data_i       ( s_soc_fll_master.data         ),
        .soc_fll_slave_ack_o        ( s_soc_fll_master.ack          ),
        .soc_fll_slave_r_data_o     ( s_soc_fll_master.r_data       ),
        .soc_fll_slave_lock_o       ( s_soc_fll_master.lock         ),

        .per_fll_slave_req_i        ( s_per_fll_master.req          ),
        .per_fll_slave_wrn_i        ( s_per_fll_master.wrn          ),
        .per_fll_slave_add_i        ( s_per_fll_master.add[1:0]     ),
        .per_fll_slave_data_i       ( s_per_fll_master.data         ),
        .per_fll_slave_ack_o        ( s_per_fll_master.ack          ),
        .per_fll_slave_r_data_o     ( s_per_fll_master.r_data       ),
        .per_fll_slave_lock_o       ( s_per_fll_master.lock         ),

        .cluster_fll_slave_req_i    ( s_cluster_fll_master.req      ),
        .cluster_fll_slave_wrn_i    ( s_cluster_fll_master.wrn      ),
        .cluster_fll_slave_add_i    ( s_cluster_fll_master.add[1:0] ),
        .cluster_fll_slave_data_i   ( s_cluster_fll_master.data     ),
        .cluster_fll_slave_ack_o    ( s_cluster_fll_master.ack      ),
        .cluster_fll_slave_r_data_o ( s_cluster_fll_master.r_data   ),
        .cluster_fll_slave_lock_o   ( s_cluster_fll_master.lock     ),

        .clk_soc_o                  ( s_soc_clk                     ),
        .clk_per_o                  ( s_periph_clk                  )
    );

    soc_interconnect_wrap #(
        .N_L2_BANKS         ( NB_L2_BANKS           ),
        .ADDR_MEM_WIDTH     ( L2_MEM_ADDR_WIDTH     ),
        .N_HWPE_PORTS       ( NB_HWPE_PORTS         ),

        .N_L2_BANKS_PRI     ( NB_L2_BANKS_PRI       ),
        .ADDR_MEM_PRI_WIDTH ( L2_MEM_ADDR_WIDTH_PRI ),

        .ROM_ADDR_WIDTH     ( ROM_ADDR_WIDTH        ),

        .AXI_32_ID_WIDTH    ( AXI_ID_OUT_WIDTH      ),
        .AXI_32_USER_WIDTH  ( AXI_USER_WIDTH        ),

        .AXI_ADDR_WIDTH     ( AXI_ADDR_WIDTH        ),
        .AXI_DATA_WIDTH     ( AXI_DATA_IN_WIDTH     ),
        .AXI_STRB_WIDTH     ( AXI_DATA_IN_WIDTH/8   ),
        .AXI_USER_WIDTH     ( AXI_USER_WIDTH        ),
        .AXI_ID_WIDTH       ( AXI_SOC_NODE_IW_OUP   )
    ) i_soc_interconnect_wrap (
        .clk_i            ( s_soc_clk           ),
        .rstn_i           ( s_soc_rstn          ),
        .test_en_i        ( dft_test_mode_i     ),
        .lint_fc_data     ( s_lint_fc_data_bus  ),
        .lint_fc_instr    ( s_lint_fc_instr_bus ),
        .lint_udma_tx     ( s_lint_udma_tx_bus  ),
        .lint_udma_rx     ( s_lint_udma_rx_bus  ),
        .lint_debug       ( s_lint_debug_bus    ),
        .lint_hwpe        ( s_lint_hwpe_bus     ),

        .axi_from_cluster ( soc_in_mst          ),
        .axi_to_cluster   ( s_data_out_bus      ),

        .apb_periph_bus   ( s_apb_periph_bus    ),
        .mem_l2_bus       ( s_mem_l2_bus        ),
        .mem_l2_pri_bus   ( s_mem_l2_pri_bus    ),
        .mem_rom_bus      ( s_mem_rom_bus       )
    );


    /* Debug Subsystem */

    dmi_jtag #(
        .IdcodeValue          ( `DMI_JTAG_IDCODE    )
    ) i_dmi_jtag (
        .clk_i                ( s_soc_clk           ),
        .rst_ni               ( s_soc_rstn          ),
        .testmode_i           ( 1'b0                ),
        .dmi_req_o            ( jtag_dmi_req        ),
        .dmi_req_valid_o      ( jtag_req_valid      ),
        .dmi_req_ready_i      ( debug_req_ready     ),
        .dmi_resp_i           ( debug_resp          ),
        .dmi_resp_ready_o     ( jtag_resp_ready     ),
        .dmi_resp_valid_i     ( jtag_resp_valid     ),
        .dmi_rst_no           (                     ), // not connected
        .tck_i                ( jtag_tck_i          ),
        .tms_i                ( jtag_tms_i          ),
        .trst_ni              ( jtag_trst_ni        ),
        .td_i                 ( jtag_tdi_i          ),
        .td_o                 ( int_td              ),
        .tdo_oe_o             (                     )
    );

   // assign hartinfo
   generate
      for(nhart_var=0;nhart_var<NrHarts;nhart_var=nhart_var+1)
        assign hartinfo[nhart_var] = '{
                                       zero1:        '0,
                                       nscratch:      2, // Debug module needs at least two scratch regs
                                       zero0:        '0,
                                       dataaccess: 1'b1, // data registers are memory mapped in the debugger
                                       datasize: dm::DataCount,
                                       dataaddr: dm::DataAddr
                                       };
   endgenerate

   generate
      for(dbg_var=0;dbg_var<NB_CORES;dbg_var=dbg_var+1)
        assign cluster_dbg_irq_valid_o[dbg_var] = dm_debug_req[CLUSTER_CORE_ID[dbg_var]];
   endgenerate

    dm_top #(
       .NrHarts           ( NrHarts                   ),
       .BusWidth          ( 32                        ),
       .SelectableHarts   ( SELECTABLE_HARTS          )
    ) i_dm_top (

       .clk_i             ( s_soc_clk                 ),
       .rst_ni            ( s_soc_rstn                ),
       .testmode_i        ( 1'b0                      ),
       .ndmreset_o        (                           ),
       .dmactive_o        (                           ), // active debug session
       .debug_req_o       ( dm_debug_req              ),
       .unavailable_i     ( ~SELECTABLE_HARTS         ),
       .hartinfo_i        ( hartinfo                  ),

       .slave_req_i       ( slave_req                 ),
       .slave_we_i        ( slave_we                  ),
       .slave_addr_i      ( slave_addr                ),
       .slave_be_i        ( slave_be                  ),
       .slave_wdata_i     ( slave_wdata               ),
       .slave_rdata_o     ( slave_rdata               ),

       .master_req_o      ( s_lint_riscv_jtag_bus.req      ),
       .master_add_o      ( s_lint_riscv_jtag_bus.add      ),
       .master_we_o       ( lint_riscv_jtag_bus_master_we  ),
       .master_wdata_o    ( s_lint_riscv_jtag_bus.wdata    ),
       .master_be_o       ( s_lint_riscv_jtag_bus.be       ),
       .master_gnt_i      ( s_lint_riscv_jtag_bus.gnt      ),
       .master_r_valid_i  ( s_lint_riscv_jtag_bus.r_valid  ),
       .master_r_rdata_i  ( s_lint_riscv_jtag_bus.r_rdata  ),

       .dmi_rst_ni        ( s_soc_rstn                ),
       .dmi_req_valid_i   ( jtag_req_valid            ),
       .dmi_req_ready_o   ( debug_req_ready           ),
       .dmi_req_i         ( jtag_dmi_req              ),
       .dmi_resp_valid_o  ( jtag_resp_valid           ),
       .dmi_resp_ready_i  ( jtag_resp_ready           ),
       .dmi_resp_o        ( debug_resp                )
    );
    assign s_lint_riscv_jtag_bus.wen = ~lint_riscv_jtag_bus_master_we;

    jtag_tap_top jtag_tap_top_i
    (
        .tck_i                    ( jtag_tck_i         ),
        .trst_ni                  ( jtag_trst_ni       ),
        .tms_i                    ( jtag_tms_i         ),
        .td_i                     ( int_td             ),
        .td_o                     ( jtag_tdo_o         ),

        .test_clk_i               ( 1'b0               ),
        .test_rstn_i              ( s_soc_rstn         ),

        .jtag_shift_dr_o          ( s_jtag_shift_dr    ),
        .jtag_update_dr_o         ( s_jtag_update_dr   ),
        .jtag_capture_dr_o        ( s_jtag_capture_dr  ),

        .axireg_sel_o             ( s_jtag_axireg_sel  ),
        .dbg_axi_scan_in_o        ( s_jtag_axireg_tdi  ),
        .dbg_axi_scan_out_i       ( s_jtag_axireg_tdo  ),
        .soc_jtag_reg_i           ( soc_jtag_reg_soc   ),
        .soc_jtag_reg_o           ( soc_jtag_reg_tap   ),
        .sel_fll_clk_o            ( s_sel_fll_clk      )
    );

    lint_jtag_wrap i_lint_jtag (
        .tck_i                    ( jtag_tck_i           ),
        .tdi_i                    ( s_jtag_axireg_tdi    ),
        .trstn_i                  ( jtag_trst_ni         ),
        .tdo_o                    ( s_jtag_axireg_tdo    ),
        .shift_dr_i               ( s_jtag_shift_dr      ),
        .pause_dr_i               ( 1'b0                 ),
        .update_dr_i              ( s_jtag_update_dr     ),
        .capture_dr_i             ( s_jtag_capture_dr    ),
        .lint_select_i            ( s_jtag_axireg_sel    ),
        .clk_i                    ( s_soc_clk            ),
        .rst_ni                   ( s_soc_rstn           ),
        .jtag_lint_master         ( s_lint_pulp_jtag_bus )
    );

    tcdm_arbiter_2x1 jtag_lint_arbiter_i
     (
        .clk_i(s_soc_clk),
        .rst_ni(s_soc_rstn),
        .tcdm_bus_1_i(s_lint_riscv_jtag_bus),
        .tcdm_bus_0_i(s_lint_pulp_jtag_bus),
        .tcdm_bus_o(s_lint_debug_bus)
    );

    apb2per #(
        .PER_ADDR_WIDTH ( 32  ),
        .APB_ADDR_WIDTH ( 32  )
    ) apb2per_newdebug_i (
        .clk_i                ( s_soc_clk               ),
        .rst_ni               ( s_soc_rstn              ),

        .PADDR                ( s_apb_debug_bus.paddr   ),
        .PWDATA               ( s_apb_debug_bus.pwdata  ),
        .PWRITE               ( s_apb_debug_bus.pwrite  ),
        .PSEL                 ( s_apb_debug_bus.psel    ),
        .PENABLE              ( s_apb_debug_bus.penable ),
        .PRDATA               ( s_apb_debug_bus.prdata  ),
        .PREADY               ( s_apb_debug_bus.pready  ),
        .PSLVERR              ( s_apb_debug_bus.pslverr ),

        .per_master_req_o     ( slave_req               ),
        .per_master_add_o     ( slave_addr              ),
        .per_master_we_o      ( slave_we                ),
        .per_master_wdata_o   ( slave_wdata             ),
        .per_master_be_o      ( slave_be                ),
        .per_master_gnt_i     ( slave_grant             ),
        .per_master_r_valid_i ( slave_valid             ),
        .per_master_r_opc_i   ( '0                      ),
        .per_master_r_rdata_i ( slave_rdata             )
     );

     assign slave_grant = slave_req;
     always_ff @(posedge s_soc_clk or negedge s_soc_rstn) begin : apb2per_valid
         if(~s_soc_rstn) begin
             slave_valid <= 0;
         end else begin
             slave_valid <= slave_grant;
         end
     end

    //********************************************************
    //*** PAD AND GPIO CONFIGURATION SIGNALS PACK ************
    //********************************************************

    generate
        for (i=0; i<32; i++) begin
            for (j=0; j<6; j++) begin
                assign gpio_cfg_o[j+6*i] = s_gpio_cfg[i][j];
            end
        end
    endgenerate

    generate
        for (i=0; i<64; i++) begin
            for (j=0; j<2; j++) begin
                assign pad_mux_o[j+2*i] = s_pad_mux[i][j];
            end
        end
    endgenerate

    generate
        for (i=0; i<64; i++) begin
            for (j=0; j<6; j++) begin
                assign pad_cfg_o[j+6*i] = s_pad_cfg[i][j];
            end
        end
    endgenerate

    //********************************************************
    //*** AXI DATA SLAVE INTERFACE UNPACK ********************
    //********************************************************

    // AXI DATA SLAVE
    assign s_data_slave.aw_writetoken  = data_slave_aw_writetoken_i  ;
    assign s_data_slave.aw_addr        = data_slave_aw_addr_i        ;
    assign s_data_slave.aw_prot        = data_slave_aw_prot_i        ;
    assign s_data_slave.aw_region      = data_slave_aw_region_i      ;
    assign s_data_slave.aw_len         = data_slave_aw_len_i         ;
    assign s_data_slave.aw_size        = data_slave_aw_size_i        ;
    assign s_data_slave.aw_burst       = data_slave_aw_burst_i       ;
     //assign s_data_slave.aw_atop        = data_slave_aw_atop_i        ;
    assign s_data_slave.aw_lock        = data_slave_aw_lock_i        ;
    assign s_data_slave.aw_cache       = data_slave_aw_cache_i       ;
    assign s_data_slave.aw_qos         = data_slave_aw_qos_i         ;
    assign s_data_slave.aw_id          = data_slave_aw_id_i          ;
    assign s_data_slave.aw_user        = data_slave_aw_user_i        ;
    assign data_slave_aw_readpointer_o = s_data_slave.aw_readpointer ;

    assign s_data_slave.ar_writetoken  = data_slave_ar_writetoken_i  ;
    assign s_data_slave.ar_addr        = data_slave_ar_addr_i        ;
    assign s_data_slave.ar_prot        = data_slave_ar_prot_i        ;
    assign s_data_slave.ar_region      = data_slave_ar_region_i      ;
    assign s_data_slave.ar_len         = data_slave_ar_len_i         ;
    assign s_data_slave.ar_size        = data_slave_ar_size_i        ;
    assign s_data_slave.ar_burst       = data_slave_ar_burst_i       ;
    assign s_data_slave.ar_lock        = data_slave_ar_lock_i        ;
    assign s_data_slave.ar_cache       = data_slave_ar_cache_i       ;
    assign s_data_slave.ar_qos         = data_slave_ar_qos_i         ;
    assign s_data_slave.ar_id          = data_slave_ar_id_i          ;
    assign s_data_slave.ar_user        = data_slave_ar_user_i        ;
    assign data_slave_ar_readpointer_o = s_data_slave.ar_readpointer ;

    assign s_data_slave.w_writetoken   = data_slave_w_writetoken_i   ;
    assign s_data_slave.w_data         = data_slave_w_data_i         ;
    assign s_data_slave.w_strb         = data_slave_w_strb_i         ;
    assign s_data_slave.w_user         = data_slave_w_user_i         ;
    assign s_data_slave.w_last         = data_slave_w_last_i         ;
    assign data_slave_w_readpointer_o  = s_data_slave.w_readpointer  ;

    assign data_slave_r_writetoken_o   = s_data_slave.r_writetoken   ;
    assign data_slave_r_data_o         = s_data_slave.r_data         ;
    assign data_slave_r_resp_o         = s_data_slave.r_resp         ;
    assign data_slave_r_last_o         = s_data_slave.r_last         ;
    assign data_slave_r_id_o           = s_data_slave.r_id           ;
    assign data_slave_r_user_o         = s_data_slave.r_user         ;
    assign s_data_slave.r_readpointer  = data_slave_r_readpointer_i  ;

    assign data_slave_b_writetoken_o   = s_data_slave.b_writetoken   ;
    assign data_slave_b_resp_o         = s_data_slave.b_resp         ;
    assign data_slave_b_id_o           = s_data_slave.b_id           ;
    assign data_slave_b_user_o         = s_data_slave.b_user         ;
    assign s_data_slave.b_readpointer  = data_slave_b_readpointer_i  ;

    //********************************************************
    //*** AXI DATA MASTER INTERFACE UNPACK *******************
    //********************************************************

    assign data_master_aw_writetoken_o  = s_data_master.aw_writetoken ;
    assign data_master_aw_addr_o        = s_data_master.aw_addr       ;
    assign data_master_aw_prot_o        = s_data_master.aw_prot       ;
    assign data_master_aw_region_o      = s_data_master.aw_region     ;
    assign data_master_aw_len_o         = s_data_master.aw_len        ;
    assign data_master_aw_size_o        = s_data_master.aw_size       ;
    //assign data_master_aw_atop_o        = s_data_master.aw_atop       ;
    assign data_master_aw_burst_o       = s_data_master.aw_burst      ;
    assign data_master_aw_lock_o        = s_data_master.aw_lock       ;
    assign data_master_aw_cache_o       = s_data_master.aw_cache      ;
    assign data_master_aw_qos_o         = s_data_master.aw_qos        ;
    assign data_master_aw_id_o          = s_data_master.aw_id         ;
    assign data_master_aw_user_o        = s_data_master.aw_user       ;
    assign s_data_master.aw_readpointer = data_master_aw_readpointer_i;

    assign data_master_ar_writetoken_o  = s_data_master.ar_writetoken ;
    assign data_master_ar_addr_o        = s_data_master.ar_addr       ;
    assign data_master_ar_prot_o        = s_data_master.ar_prot       ;
    assign data_master_ar_region_o      = s_data_master.ar_region     ;
    assign data_master_ar_len_o         = s_data_master.ar_len        ;
    assign data_master_ar_size_o        = s_data_master.ar_size       ;
    assign data_master_ar_burst_o       = s_data_master.ar_burst      ;
    assign data_master_ar_lock_o        = s_data_master.ar_lock       ;
    assign data_master_ar_cache_o       = s_data_master.ar_cache      ;
    assign data_master_ar_qos_o         = s_data_master.ar_qos        ;
    assign data_master_ar_id_o          = s_data_master.ar_id         ;
    assign data_master_ar_user_o        = s_data_master.ar_user       ;
    assign s_data_master.ar_readpointer = data_master_ar_readpointer_i;

    assign data_master_w_writetoken_o   = s_data_master.w_writetoken  ;
    assign data_master_w_data_o         = s_data_master.w_data        ;
    assign data_master_w_strb_o         = s_data_master.w_strb        ;
    assign data_master_w_user_o         = s_data_master.w_user        ;
    assign data_master_w_last_o         = s_data_master.w_last        ;
    assign s_data_master.w_readpointer  = data_master_w_readpointer_i ;

    assign s_data_master.r_writetoken   = data_master_r_writetoken_i  ;
    assign s_data_master.r_data         = data_master_r_data_i        ;
    assign s_data_master.r_resp         = data_master_r_resp_i        ;
    assign s_data_master.r_last         = data_master_r_last_i        ;
    assign s_data_master.r_id           = data_master_r_id_i          ;
    assign s_data_master.r_user         = data_master_r_user_i        ;
    assign data_master_r_readpointer_o  = s_data_master.r_readpointer ;

    assign s_data_master.b_writetoken   = data_master_b_writetoken_i  ;
    assign s_data_master.b_resp         = data_master_b_resp_i        ;
    assign s_data_master.b_id           = data_master_b_id_i          ;
    assign s_data_master.b_user         = data_master_b_user_i        ;
    assign data_master_b_readpointer_o  = s_data_master.b_readpointer ;

endmodule

// Local Variables:
// verilog-indent-level: 4
// verilog-indent-level-module: 4
// verilog-indent-level-declaration: 4
// verilog-indent-level-behavioral: 4
// verilog-case-indent: 4
// verilog-cexp-indent: 4
// End:
