// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

`include "pulp_soc_defines.sv"

`ifndef PULP_FPGA_EMUL
 `ifdef SYNTHESIS
  `define ASIC_SYNTHESIS
 `endif
`endif

module fc_subsystem #(
    parameter CORE_TYPE           = 0,
    parameter PULP_XPULP          = 1,
    parameter USE_FPU             = 1,
    parameter ZFINX               = 0,
    parameter USE_HWPE            = 1,
    parameter EVENT_ID_WIDTH      = 8,
    parameter PER_ID_WIDTH        = 32,
    parameter NB_HWPE_PORTS       = 4,
    parameter PULP_SECURE         = 1,
    parameter TB_RISCV            = 0,
    parameter CORE_ID             = 4'h0,
    parameter CLUSTER_ID          = 6'h1F
) (
    input  logic                      clk_i,
    input  logic                      rst_ni,
    input  logic                      test_en_i,

    input logic           wdt_reset_i,

    XBAR_TCDM_BUS.Master              l2_data_master,
    XBAR_TCDM_BUS.Master              l2_instr_master,
    XBAR_TCDM_BUS.Master              l2_hwpe_master [NB_HWPE_PORTS-1:0],
    APB_BUS.Slave                     apb_slave_eu,
    APB_BUS.Slave                     apb_slave_hwpe,

    input  logic                      fetch_en_i,
    input  logic [31:0]               boot_addr_i,
    input  logic                      debug_req_i,

    input  logic                      event_fifo_valid_i,
    output logic                      event_fifo_fulln_o,
    input  logic [EVENT_ID_WIDTH-1:0] event_fifo_data_i, // goes indirectly to core interrupt
    input  logic [31:0]               events_i, // goes directly to core interrupt, should be called irqs

    input  logic                      plic_irq_valid_i,
    output logic                      plic_irq_ready_o,

    output logic [1:0]                hwpe_events_o,

    output logic                      supervisor_mode_o
);

    import cv32e40p_apu_core_pkg::*;

    // Number of performance counters. As previously in RI5CY (riscv_cs_registers.sv),
    // we distinguish between:
    // (a) ASIC implementation: 1 performance counter active
    // (b) RTL simulation/FPGA emulation: 16 performance counters active, one for each event

    `ifdef ASIC_SYNTHESIS
      localparam int unsigned NUM_MHPMCOUNTERS = 1;
    `else
      localparam int unsigned NUM_MHPMCOUNTERS = 16;
    `endif

    // Interrupt signals
    logic        core_irq_req   ;
    logic        core_irq_sec   ;
    logic [4:0]  core_irq_id    ;
    logic [4:0]  core_irq_ack_id;
    logic        core_irq_ack   ;
    logic [14:0] core_irq_fast  ;
    logic [31:0] core_irq_x     ;

    logic [3:0]  irq_ack_id;

    // Signals for OBI-PULP conversion
    logic        obi_instr_req;
    logic        pulp_instr_req;

    // Boot address, core id, cluster id, fethc enable and core_status
    logic [31:0] boot_addr        ;
    logic        fetch_en_int     ;
    logic        core_busy_int    ;
    logic        perf_counters_int;
    logic [31:0] hart_id;

    //EU signals
    logic core_clock_en;
    logic fetch_en_eu  ;

    //Core Instr Bus
    logic [31:0] core_instr_addr, core_instr_rdata;
    logic        core_instr_req, core_instr_gnt, core_instr_rvalid, core_instr_err;

    //Core Data Bus
    logic [31:0] core_data_addr, core_data_rdata, core_data_wdata;
    logic        core_data_req, core_data_gnt, core_data_rvalid;
    logic        core_data_we  ;
    logic [ 3:0]  core_data_be ;
    logic is_scm_instr_req, is_scm_data_req;

    logic core_rst;

    assign perf_counters_int = 1'b0;
    assign fetch_en_int      = fetch_en_eu & fetch_en_i;

    assign hart_id = {21'b0, CLUSTER_ID[5:0], 1'b0, CORE_ID[3:0]};

    XBAR_TCDM_BUS core_data_bus ();
    XBAR_TCDM_BUS core_instr_bus ();

    // APU Core to FP Wrapper
    logic                               apu_req;
    logic [    APU_NARGS_CPU-1:0][31:0] apu_operands;
    logic [      APU_WOP_CPU-1:0]       apu_op;
    logic [ APU_NDSFLAGS_CPU-1:0]       apu_flags;


    // APU FP Wrapper to Core
    logic                               apu_gnt;
    logic                               apu_rvalid;
    logic [                 31:0]       apu_rdata;
    logic [ APU_NUSFLAGS_CPU-1:0]       apu_rflags;

    //********************************************************
    //************ CORE DEMUX (TCDM vs L2) *******************
    //********************************************************
    assign l2_data_master.req    = core_data_req;
    assign l2_data_master.add    = core_data_addr;
    assign l2_data_master.wen    = ~core_data_we;
    assign l2_data_master.wdata  = core_data_wdata;
    assign l2_data_master.be     = core_data_be;
    assign core_data_gnt         = l2_data_master.gnt;
    assign core_data_rvalid      = l2_data_master.r_valid;
    assign core_data_rdata       = l2_data_master.r_rdata;
    assign core_data_err         = l2_data_master.r_opc;


    assign l2_instr_master.req   = core_instr_req;
    assign l2_instr_master.add   = core_instr_addr;
    assign l2_instr_master.wen   = 1'b1;
    assign l2_instr_master.wdata = '0;
    assign l2_instr_master.be    = 4'b1111;
    assign core_instr_gnt        = l2_instr_master.gnt;
    assign core_instr_rvalid     = l2_instr_master.r_valid;
    assign core_instr_rdata      = l2_instr_master.r_rdata;
    assign core_instr_err        = l2_instr_master.r_opc;

    //********************************************************
    //************ RISCV CORE ********************************
    //********************************************************
    assign core_rst = rst_ni  & ~wdt_reset_i;

    assign boot_addr = boot_addr_i;
`ifndef PULP_FPGA_EMUL
  `ifdef SYNTHESIS
    cv32e40p_core #(
  `else
    cv32e40p_wrapper #(
  `endif
`else
    cv32e40p_core #(
`endif
        .PULP_XPULP       (PULP_XPULP),
        .PULP_CLUSTER     (0),
        .FPU              (USE_FPU),
        .PULP_ZFINX       (ZFINX),
        .NUM_MHPMCOUNTERS (NUM_MHPMCOUNTERS)
    ) FC_CORE_i (

        // Clock and Reset
        .clk_i                (clk_i),
        .rst_ni               (rst_ni),

        // Core ID, Cluster ID, debug mode halt address and boot address are considered more or less static
        .pulp_clock_en_i      (clock_en_i ),
        .scan_cg_en_i         (test_mode_i),
        .boot_addr_i          (boot_addr),
        .mtvec_addr_i         (),
        .dm_halt_addr_i       (32'h1A110800),
        .hart_id_i            (hart_id),
        .dm_exception_addr_i  (32'h1A11080c),

        // Instruction memory interface
        .instr_req_o           (obi_instr_req),
        .instr_gnt_i           (core_instr_gnt),
        .instr_rvalid_i        (core_instr_rvalid),
        .instr_addr_o          (core_instr_addr),
        .instr_rdata_i         (core_instr_rdata),

        // Data memory interface
        .data_req_o            (core_data_req),
        .data_gnt_i            (core_data_gnt),
        .data_rvalid_i         (core_data_rvalid),
        .data_we_o             (core_data_we),
        .data_be_o             (core_data_be),
        .data_addr_o           (core_data_addr),
        .data_wdata_o          (core_data_wdata),
        .data_rdata_i          (core_data_rdata),

        // apu-interconnect
        // handshake signals
        .apu_req_o             (apu_req),
        .apu_gnt_i             (apu_gnt),
        // request channel
        .apu_operands_o        (apu_operands),
        .apu_op_o              (apu_op),
        .apu_flags_o           (apu_flags),
        // response channel
        .apu_rvalid_i          (apu_rvalid),
        .apu_result_i          (apu_rdata),
        .apu_flags_i           (apu_rflags),

        // Interrupt inputs
        .irq_i                 (core_irq_x),  // CLINT interrupts + CLINT extension interrupts
        .irq_ack_o             (core_irq_ack),
        .irq_id_o              (core_irq_ack_id),

        // Debug Interface
        .debug_req_i           (debug_req_i),
        .debug_havereset_o     (),
        .debug_running_o       (),
        .debug_halted_o        (),

        // CPU Control Signals
        .fetch_enable_i        (fetch_en_int),
        .core_sleep_o          ()
    );

    // OBI-PULP adapter
    obi_pulp_adapter i_obi_pulp_adapter (
        .rst_ni       (rst_ni),
        .clk_i        (clk_i),
        .core_req_i   (obi_instr_req),
        .mem_gnt_i    (core_instr_gnt),
        .mem_rvalid_i (core_instr_rvalid),
        .mem_req_o    (pulp_instr_req)
      );
    assign core_instr_req = pulp_instr_req;

    assign supervisor_mode_o = 1'b1;

    //// remap ack ID for SoC Event FIFO
    //always_comb begin : gen_core_irq_ack_id
    //    if (irq_ack_id == 10) begin
    //        core_irq_ack_id = 26;
    //    end else begin
    //        core_irq_ack_id = {1'b0, irq_ack_id};
    //    end
    //end

    always_comb begin : gen_core_irq_x
        core_irq_x = '0;
        if (core_irq_req) begin
            core_irq_x[core_irq_id] = 1'b1;
        end
    end

    apb_interrupt_cntrl #(.PER_ID_WIDTH(PER_ID_WIDTH)) fc_eu_i (
        .clk_i              ( clk_i              ),
        .rst_ni             ( rst_ni             ),
        .test_mode_i        ( test_en_i          ),
        .events_i           ( events_i           ),
        .event_fifo_valid_i ( event_fifo_valid_i ),
        .event_fifo_fulln_o ( event_fifo_fulln_o ),
        .event_fifo_data_i  ( event_fifo_data_i  ),
        .plic_irq_valid_i,
        .plic_irq_ready_o,
        .core_secure_mode_i ( 1'b0               ),
        .core_irq_id_o      ( core_irq_id        ),
        .core_irq_req_o     ( core_irq_req       ),
        .core_irq_ack_i     ( core_irq_ack       ),
        .core_irq_id_i      ( core_irq_ack_id    ),
        .core_irq_sec_o     ( /* SECURE IRQ */   ),
        .core_clock_en_o    ( core_clock_en      ),
        .fetch_en_o         ( fetch_en_eu        ),
        .apb_slave          ( apb_slave_eu       )
    );


    generate
    if(USE_HWPE) begin : fc_hwpe_gen
        fc_hwpe #(
            .N_MASTER_PORT ( NB_HWPE_PORTS ),
            .ID_WIDTH      ( 2             )
        ) i_fc_hwpe (
            .clk_i             ( clk_i          ),
            .rst_ni            ( rst_ni         ),
            .test_mode_i       ( test_en_i      ),
            .hwacc_xbar_master ( l2_hwpe_master ),
            .hwacc_cfg_slave   ( apb_slave_hwpe ),
            .evt_o             ( hwpe_events_o  ),
            .busy_o            (                )
        );
    end
    else begin : no_fc_hwpe_gen
        assign hwpe_events_o = '0;
        assign apb_slave_hwpe.prdata  = '0;
        assign apb_slave_hwpe.pready  = '0;
        assign apb_slave_hwpe.pslverr = '0;
        for(genvar ii=0; ii<NB_HWPE_PORTS; ii++) begin
            assign l2_hwpe_master[ii].req   = '0;
            assign l2_hwpe_master[ii].wen   = '0;
            assign l2_hwpe_master[ii].wdata = '0;
            assign l2_hwpe_master[ii].be    = '0;
            assign l2_hwpe_master[ii].add   = '0;
        end
    end
    endgenerate


    //*************************************
    //****** APU INTERFACE WITH FPU *******
    //*************************************

`ifdef FPU_SOC
    cv32e40p_fp_wrapper #(
        .FP_DIVSQRT (1)
    ) fp_wrapper_i (
        .clk_i         (clk_i),
        .rst_ni        (rst_ni),
        .apu_req_i     (apu_req),
        .apu_gnt_o     (apu_gnt),
        .apu_operands_i(apu_operands),
        .apu_op_i      (apu_op),
        .apu_flags_i   (apu_flags),
        .apu_rvalid_o  (apu_rvalid),
        .apu_rdata_o   (apu_rdata),
        .apu_rflags_o  (apu_rflags)
    );
`else
    assign apu_req      = 1'b0;
    assign apu_gnt      = 1'b0;
    assign apu_operands = 1'b0;
    assign apu_op       = 1'b0;
    assign apu_flags    = 1'b0;
    assign apu_rvalid   = 1'b0;
    assign apu_rdata    = 1'b0;
    assign apu_rflags   = 1'b0;
`endif // !`ifdef FPU_SOC

endmodule
