// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.


`include "pulp_soc_defines.sv"
`include "axi/typedef.svh"
`include "axi/assign.svh"

module pulp_soc import dm::*; #(
    parameter CORE_TYPE          = 0,
    parameter PULP_XPULP         = 1,
    parameter USE_FPU            = 1,
    parameter USE_HWPE           = 1,
    parameter USE_CLUSTER_EVENT  = 1,
    parameter ZFINX              = 0,
    parameter N_PERF_COUNTERS    = 1,
    parameter SIM_STDOUT         = 1,
    parameter AXI_ADDR_WIDTH     = 32,
    parameter AXI_DATA_IN_WIDTH  = 64,
    parameter AXI_DATA_OUT_S2C_WIDTH = 32,
    parameter AXI_DATA_OUT_S2E_WIDTH = 64,
    parameter AXI_ID_IN_WIDTH    = 7,
    parameter AXI_ID_OUT_S2C_WIDTH = 5,
    parameter AXI_ID_OUT_S2E_WIDTH = 6,
    parameter AXI_USER_WIDTH     = 6,
    parameter AXI_STRB_WIDTH_IN  = AXI_DATA_IN_WIDTH/8,
    parameter AXI_STRB_WIDTH_S2C_OUT = AXI_DATA_OUT_S2C_WIDTH/8,
    parameter AXI_STRB_WIDTH_S2E_OUT = AXI_DATA_OUT_S2E_WIDTH/8,
    parameter BUFFER_WIDTH       = 8,
    parameter C2S_AW_WIDTH       = 80,
    parameter C2S_W_WIDTH        = 79,
    parameter C2S_B_WIDTH        = 15,
    parameter C2S_AR_WIDTH       = 74,
    parameter C2S_R_WIDTH        = 80,
    parameter S2C_AW_WIDTH       = 78,
    parameter S2C_W_WIDTH        = 43,
    parameter S2C_B_WIDTH        = 13,
    parameter S2C_AR_WIDTH       = 72,
    parameter S2C_R_WIDTH        = 46,
    parameter LOG_DEPTH          = 3,
    parameter EVNT_WIDTH         = 8,
    parameter NB_CORES           = 8,
    parameter NB_HWPE_PORTS      = 4,
    parameter NGPIO              = 32,
    parameter NBIT_PADCFG        = 4, //Must not be changed as other parts
                                      //downstreams are not parametrci

    parameter int unsigned N_UART = 1,
    parameter int unsigned N_SPI  = 1,
    parameter int unsigned N_I2C  = 2,
    parameter int unsigned N_I2C_SLV  = 2,

    parameter int unsigned N_L2_BANKS = 0,
    parameter int unsigned N_L2_BANKS_PRI = 0,
    parameter int unsigned L2_BANK_SIZE = 0,
    parameter int unsigned L2_BANK_SIZE_PRI = 0,
    parameter int unsigned L2_SIZE = 0,
    parameter int unsigned NUM_INTERRUPTS = 0,
    parameter int unsigned MACRO_ROM = 0,
    parameter int unsigned USE_CLUSTER = 1
) (
    input  logic                          soc_clk_i,
    input  logic                          periph_clk_i,
    input  logic                          ref_clk_i,
    input  logic                          test_clk_i,
    input  logic                          soc_rst_ni,
    input  logic                          cluster_rst_ni,

    input  logic                          dft_test_mode_i,
    input  logic                          dft_cg_enable_i,
    input  logic                          mode_select_i,
    input  logic                          bootsel_valid_i,
    input  logic [2:0]                    bootsel_i,

    input  logic                          fc_fetch_en_valid_i,
    input  logic                          fc_fetch_en_i,

    // AXI interfaces to outside of control pulp
    AXI_BUS.Slave                         axi_ext_slv,  // from ext
    AXI_BUS.Master                        axi_ext_mst,

    // TCDM interfaces to memory cuts (all are placed outside of control-pulp)
    XBAR_TCDM_BUS.Master                  s_mem_l2_bus[N_L2_BANKS],
    XBAR_TCDM_BUS.Master                  s_mem_l2_pri_bus[N_L2_BANKS_PRI],

    // APB interfaces to configure external IPs
    APB_BUS.Master                        apb_clk_ctrl_bus,
    output logic                          clk_mux_sel_o,
    APB_BUS.Master                        apb_serial_link_bus,
    APB_BUS.Master                        apb_pad_cfg_bus,

    output logic                          cluster_fetch_enable_o,
    output logic [63:0]                   cluster_boot_addr_o,
    output logic                          cluster_test_en_o,
    output logic                          cluster_pow_o,
    output logic                          cluster_byp_o,
    output logic                          cluster_rst_reg_no,
    output logic                          cluster_irq_o,

    // AXI4 SLAVE
    input logic [LOG_DEPTH:0]                         async_data_slave_aw_wptr_i,
    input logic [2**LOG_DEPTH-1:0][C2S_AW_WIDTH-1:0]  async_data_slave_aw_data_i,
    output logic [LOG_DEPTH:0]                        async_data_slave_aw_rptr_o,

    // READ ADDRESS CHANNEL
    input logic [LOG_DEPTH:0]                         async_data_slave_ar_wptr_i,
    input logic [2**LOG_DEPTH-1:0][C2S_AR_WIDTH-1:0]  async_data_slave_ar_data_i,
    output logic [LOG_DEPTH:0]                        async_data_slave_ar_rptr_o,

    // WRITE DATA CHANNEL
    input logic [LOG_DEPTH:0]                         async_data_slave_w_wptr_i,
    input logic [2**LOG_DEPTH-1:0][C2S_W_WIDTH-1:0]   async_data_slave_w_data_i,
    output logic [LOG_DEPTH:0]                        async_data_slave_w_rptr_o,

    // READ DATA CHANNEL
    output logic [LOG_DEPTH:0]                        async_data_slave_r_wptr_o,
    output logic [2**LOG_DEPTH-1:0][C2S_R_WIDTH-1:0]  async_data_slave_r_data_o,
    input logic [LOG_DEPTH:0]                         async_data_slave_r_rptr_i,

    // WRITE RESPONSE CHANNEL
    output logic [LOG_DEPTH:0]                        async_data_slave_b_wptr_o,
    output logic [2**LOG_DEPTH-1:0][C2S_B_WIDTH-1:0]  async_data_slave_b_data_o,
    input logic [LOG_DEPTH:0]                         async_data_slave_b_rptr_i,

    // AXI4 MASTER
    output logic [LOG_DEPTH:0]                        async_data_master_aw_wptr_o,
    output logic [2**LOG_DEPTH-1:0][S2C_AW_WIDTH-1:0] async_data_master_aw_data_o,
    input logic [LOG_DEPTH:0]                         async_data_master_aw_rptr_i,

    // READ ADDRESS CHANNEL
    output logic [LOG_DEPTH:0]                        async_data_master_ar_wptr_o,
    output logic [2**LOG_DEPTH-1:0][S2C_AR_WIDTH-1:0] async_data_master_ar_data_o,
    input logic [LOG_DEPTH:0]                         async_data_master_ar_rptr_i,

    // WRITE DATA CHANNEL
    output logic [LOG_DEPTH:0]                        async_data_master_w_wptr_o,
    output logic [2**LOG_DEPTH-1:0][S2C_W_WIDTH-1:0]  async_data_master_w_data_o,
    input logic [LOG_DEPTH:0]                         async_data_master_w_rptr_i,

    // READ DATA CHANNEL
    input logic [LOG_DEPTH:0]                         async_data_master_r_wptr_i,
    input logic [2**LOG_DEPTH-1:0][S2C_R_WIDTH-1:0]   async_data_master_r_data_i,
    output logic [LOG_DEPTH:0]                        async_data_master_r_rptr_o,

    // WRITE RESPONSE CHANNEL
    input logic [LOG_DEPTH:0]                         async_data_master_b_wptr_i,
    input logic [2**LOG_DEPTH-1:0][S2C_B_WIDTH-1:0]   async_data_master_b_data_i,
    output logic [LOG_DEPTH:0]                        async_data_master_b_rptr_o,

    output logic [BUFFER_WIDTH-1:0]                   cluster_events_wt_o,
    input logic [BUFFER_WIDTH-1:0]                    cluster_events_rp_i,
    output logic [EVNT_WIDTH-1:0]                     cluster_events_da_o,
    input logic                                       cluster_busy_i,
    output logic                                      dma_pe_evt_ack_o,
    input logic                                       dma_pe_evt_valid_i,
    output logic                                      dma_pe_irq_ack_o,
    input logic                                       dma_pe_irq_valid_i,
    output logic                                      pf_evt_ack_o,
    input logic                                       pf_evt_valid_i,
    ///////////////////////////////////////////////////
    //      To I/O Controller and padframe           //
    ///////////////////////////////////////////////////

    input  logic [NGPIO-1:0]                  gpio_in_i,
    output logic [NGPIO-1:0]                  gpio_out_o,
    output logic [NGPIO-1:0]                  gpio_dir_o,
    output logic [NGPIO-1:0][NBIT_PADCFG-1:0] gpio_cfg_o,

    output logic [N_UART-1:0]             uart_tx_o,
    input  logic [N_UART-1:0]             uart_rx_i,
    output logic [3:0]                    timer_ch0_o,
    output logic [3:0]                    timer_ch1_o,
    output logic [3:0]                    timer_ch2_o,
    output logic [3:0]                    timer_ch3_o,

    input  logic [N_I2C-1:0]              i2c_scl_i,
    output logic [N_I2C-1:0]              i2c_scl_o,
    output logic [N_I2C-1:0]              i2c_scl_oe_o,
    input  logic [N_I2C-1:0]              i2c_sda_i,
    output logic [N_I2C-1:0]              i2c_sda_o,
    output logic [N_I2C-1:0]              i2c_sda_oe_o,

    input logic  [N_I2C_SLV-1:0]          i2c_slv_scl_i,
    output logic [N_I2C_SLV-1:0]          i2c_slv_scl_o,
    output logic [N_I2C_SLV-1:0]          i2c_slv_scl_oe_o,
    input logic  [N_I2C_SLV-1:0]          i2c_slv_sda_i,
    output logic [N_I2C_SLV-1:0]          i2c_slv_sda_o,
    output logic [N_I2C_SLV-1:0]          i2c_slv_sda_oe_o,

    output logic [N_SPI-1:0]              spi_clk_o,
    output logic [N_SPI-1:0][3:0]         spi_csn_o,
    output logic [N_SPI-1:0][3:0]         spi_oen_o,
    output logic [N_SPI-1:0][3:0]         spi_sdo_o,
    input  logic [N_SPI-1:0][3:0]         spi_sdi_i,

    input  logic                          spi_clk_i,
    input  logic                          spi_csn_i,
    output logic [3:0]                    spi_oen_slv_o,
    output logic [3:0]                    spi_sdo_slv_o,
    input  logic [3:0]                    spi_sdi_slv_i,

    //inter-socket mux signal
    output logic                          sel_spi_dir_o,
    output logic                          sel_i2c_mux_o,

    // jtag debug
    input logic                          jtag_tck_i,
    input logic                          jtag_trst_ni,
    input logic                          jtag_tms_i,
    input logic                          jtag_tdi_i,
    output logic                         jtag_tdo_o,
    output logic [NB_CORES-1:0]          cluster_dbg_irq_valid_o,

    // watch dog timer alarm
    output logic [1:0]                    wdt_alert_o,
    input  logic                          wdt_alert_clear_i,

    // external interrupts
    input logic                           scg_irq_i,
    input logic                           scp_irq_i,
    input logic                           scp_secure_irq_i,
    input logic [71:0]                    mbox_irq_i,
    input logic [71:0]                    mbox_secure_irq_i
);

    localparam int unsigned AXI_DATA_EXT_WIDTH = 64;

    localparam int unsigned CLK_CTRL_ADDR_WIDTH = 32;
    localparam int unsigned CLK_CTRL_DATA_WIDTH = 32;

    localparam L2_MEM_ADDR_WIDTH     = $clog2(L2_BANK_SIZE * N_L2_BANKS) - $clog2(N_L2_BANKS);    // 2**L2_MEM_ADDR_WIDTH rows (64bit each) in L2 --> TOTAL L2 SIZE = 8byte * 2^L2_MEM_ADDR_WIDTH

    localparam ROM_ADDR_WIDTH        = 13;

    localparam FC_CORE_CLUSTER_ID    = 6'd31;
    localparam CL_CORE_CLUSTER_ID    = 6'd0;

    localparam FC_CORE_CORE_ID       = 4'd0;
    localparam FC_CORE_MHARTID       = {FC_CORE_CLUSTER_ID, 1'b0, FC_CORE_CORE_ID};

    //  PULP RISC-V cores have not continguos MHARTID.
    //  This leads to set the number of HARTS >= the maximum value of the MHARTID.
    //  In this case, the MHARD ID is {FC_CORE_CLUSTER_ID,1'b0,FC_CORE_CORE_ID} --> 996 (1024 chosen as power of 2)
    //  To avoid paying 1024 flip flop for each number of harts's related register, we implemented
    //  the masking parameter, aka SELECTABLE_HARTS.
    //  In One-Hot-Encoding way, you select 1 when that MHARTID-related HART can actally be selected.
    //  e.g. if you have 2 core with MHART 10 and 5, you select NrHarts=16 and SELECTABLE_HARTS = (1<<10) | (1<<5).
    //  This mask will be used to generated only the flip flop needed and the constant-propagator engine of the synthesizer
    //  will remove the other flip flops and related logic.

    localparam NrHarts                               = 1024;

    // this is a constant expression
    function logic [NrHarts-1:0] SEL_HARTS_FX();
        SEL_HARTS_FX = (1 << FC_CORE_MHARTID);
        for (int i = 0; i < NB_CORES; i++) begin
            SEL_HARTS_FX |= (1 << {CL_CORE_CLUSTER_ID, 1'b0, i[3:0]});
        end
    endfunction

    // Each hart with hartid=x sets the x'th bit in SELECTABLE_HARTS
    localparam logic [NrHarts-1:0] SELECTABLE_HARTS = SEL_HARTS_FX();

    // cluster core ids gathere as vector for convenience
    logic [NB_CORES-1:0][10:0] cluster_core_id;
    for (genvar i = 0; i < NB_CORES; i++) begin : gen_cluster_core_id
        assign cluster_core_id[i] = {CL_CORE_CLUSTER_ID, 1'b0, i[3:0]};
    end

    localparam dm::hartinfo_t RI5CY_HARTINFO = '{
       zero1:        '0,
       nscratch:      2, // Debug module needs at least two scratch regs
       zero0:        '0,
       dataaccess: 1'b1, // data registers are memory mapped in the debugger
       datasize: dm::DataCount,
       dataaddr: dm::DataAddr
    };

    dm::hartinfo_t [NrHarts-1:0] hartinfo;

    /*
       This module has been tested only with the default parameters.
    */

    //********************************************************
    //***************** SIGNALS DECLARATION ******************
    //********************************************************
    logic [ 1:0]           s_fc_hwpe_events;
    logic [31:0]           s_fc_events;

    logic [7:0]            s_soc_events_ack;
    logic [7:0]            s_soc_events_val;

    logic                  s_timer_lo_event;
    logic                  s_timer_hi_event;

    logic [EVNT_WIDTH-1:0] s_cl_event_data ;
    logic                  s_cl_event_valid;
    logic                  s_cl_event_ready;

    logic [EVNT_WIDTH-1:0] s_fc_event_data ;
    logic                  s_fc_event_valid;
    logic                  s_fc_event_ready;

    logic [7:0][31:0]      s_apb_mpu_rules;
    logic                  s_supervisor_mode;

    logic [31:0]           s_fc_bootaddr;

    logic                  s_periph_clk;
    logic                  s_soc_clk;
    logic                  s_soc_rstn;
    logic                  s_cluster_rstn;
    logic                  s_sel_clk;

    logic                  s_dma_pe_evt;
    logic                  s_dma_pe_irq;
    logic                  s_pf_evt;

    logic                  s_fc_fetchen;
    logic [NrHarts-1:0]    dm_debug_req;

    logic                  jtag_req_valid;
    logic                  debug_req_ready;
    logic                  jtag_resp_ready;
    logic                  jtag_resp_valid;
    dm::dmi_req_t          jtag_dmi_req;
    dm::dmi_resp_t         debug_resp;
    logic                  slave_grant, slave_valid, slave_req , slave_we;
    logic                  [31:0] slave_addr, slave_wdata, slave_rdata;
    logic                  [3:0]  slave_be;
    logic                  lint_riscv_jtag_bus_master_we;
    logic                  int_td;

    logic                  master_req;
    logic [31:0]           master_add;
    logic                  master_we;
    logic [31:0]           master_wdata;
    logic [3:0]            master_be;
    logic                  master_gnt;
    logic                  master_r_valid;
    logic [31:0]           master_r_rdata;


    logic [7:0]            soc_jtag_reg_tap;
    logic [7:0]            soc_jtag_reg_soc;


    logic                  spi_master0_csn3, spi_master0_csn2;

    // sdma
    logic s_sdma_term_event, s_sdma_busy;


    // tap to lint wrap
    logic                  s_jtag_shift_dr;
    logic                  s_jtag_update_dr;
    logic                  s_jtag_capture_dr;
    logic                  s_jtag_axireg_sel;
    logic                  s_jtag_axireg_tdi;
    logic                  s_jtag_axireg_tdo;

    APB_BUS                s_apb_eu_bus ();
    APB_BUS                s_apb_clic_bus ();
    APB_BUS                s_apb_hwpe_bus ();
    APB_BUS                s_apb_debug_bus();
    APB_BUS                s_apb_sdma_bus();

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH ), //64
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_data_in_bus (); // from cluster

     AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH ), //64
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_axi_tcdm_sdma_mst (); // to/from tcdm through sensor dma

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_S2C_WIDTH), //32
        .AXI_ID_WIDTH   ( AXI_ID_OUT_S2C_WIDTH  ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_data_out_bus (); // to cluster

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_S2C_WIDTH), //32
        .AXI_ID_WIDTH   ( AXI_ID_OUT_S2C_WIDTH  ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_axi_ext_core_mst (); // to ext from FC core
 
    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_S2E_WIDTH), //64
        .AXI_ID_WIDTH   ( AXI_ID_OUT_S2E_WIDTH  ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_axi_ext_core_dw_mst (); // to ext from FC core

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_S2E_WIDTH), //64
        .AXI_ID_WIDTH   ( AXI_ID_OUT_S2E_WIDTH  ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
    ) s_axi_ext_sdma_mst (); // to/from ext from sensor DMA

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( AXI_DATA_OUT_S2E_WIDTH ), //64
        .AXI_ID_WIDTH   ( AXI_ID_OUT_S2E_WIDTH   ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     )
    ) axi_mux_ext_slv[2]();
    // Wrap FC core and sdma interfaces to an array of interfaces
    `AXI_ASSIGN(axi_mux_ext_slv[0], s_axi_ext_core_dw_mst) // FC core
    `AXI_ASSIGN(axi_mux_ext_slv[1], s_axi_ext_sdma_mst) // sdma
    
    ////////////////////
    // AXI Mux inputs //
    ////////////////////

    // Route cluster/ext to 1 Mux
    localparam int unsigned N_EXT_MASTERS_TO_SOC = 3; //cl, ext, sdma

    // Route i2c slvs and spi slv to 1 Mux
    localparam int unsigned N_EXT_MASTERS_TO_SOC_PERIPH = 3; // spi_slv, i2c_slv_1, i2c_slv_2

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( 32 ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH    ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     )
    ) s_axi_spi (); // from spi_slv

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( 32 ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH    ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     )
    ) axi_i2c_slv_bmc (); // from i2c_slv_1

    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( 32 ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH    ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     )
    ) axi_i2c_slv_1 (); // from i2c_slv_2

    // Wrap into single interface
    AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( AXI_DATA_IN_WIDTH  ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH    ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     )
    ) ext_masters_to_soc [N_EXT_MASTERS_TO_SOC-1:0] ();

     AXI_BUS #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH     ),
        .AXI_DATA_WIDTH ( 32 ),
        .AXI_ID_WIDTH   ( AXI_ID_IN_WIDTH    ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH     )
    ) ext_masters_to_soc_periph [N_EXT_MASTERS_TO_SOC_PERIPH-1:0] ();

    // axi_a32_d64
    `AXI_ASSIGN(ext_masters_to_soc[0], s_data_in_bus);    // from cluster
    `AXI_ASSIGN(ext_masters_to_soc[1], axi_ext_slv);      // from ext
    `AXI_ASSIGN(ext_masters_to_soc[2], s_axi_tcdm_sdma_mst); // from sdma

    // axi_a32_d32
    `AXI_ASSIGN(ext_masters_to_soc_periph[0], s_axi_spi);        // from spi_slv
    `AXI_ASSIGN(ext_masters_to_soc_periph[1], axi_i2c_slv_1);    // from i2c_slv_1
    `AXI_ASSIGN(ext_masters_to_soc_periph[2], axi_i2c_slv_bmc);  // from i2c_slv_2

    //assign s_data_out_bus.aw_atop = 6'b0;

    APB_BUS s_apb_periph_bus ();

    XBAR_TCDM_BUS s_mem_rom_bus ();

    XBAR_TCDM_BUS s_lint_debug_bus();
    XBAR_TCDM_BUS s_lint_pulp_jtag_bus();
    XBAR_TCDM_BUS s_lint_riscv_jtag_bus();
    XBAR_TCDM_BUS s_lint_udma_tx_bus ();
    XBAR_TCDM_BUS s_lint_udma_rx_bus ();
    XBAR_TCDM_BUS s_lint_fc_data_bus ();
    XBAR_TCDM_BUS s_lint_fc_instr_bus ();
    XBAR_TCDM_BUS s_lint_fc_shadow_bus ();
    XBAR_TCDM_BUS s_lint_hwpe_bus[NB_HWPE_PORTS]();

    `ifdef REMAP_ADDRESS
        logic [3:0] base_addr_int;
        assign base_addr_int = 4'b0001; //FIXME attach this signal somewhere in the soc peripherals --> IGOR
    `endif

   // Feed FC domain with soc_clk
   assign s_soc_clk = soc_clk_i;
   assign clk_mux_sel_o = s_sel_clk;
   // Feed FC domain with soc_rst_ni
   assign s_soc_rstn = soc_rst_ni;

   // If you want to connect a real PULP cluster you also need a cluster_busy_i signal

   `AXI_TYPEDEF_AW_CHAN_T(c2s_aw_chan_t,logic[AXI_ADDR_WIDTH-1:0],logic[AXI_ID_IN_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_W_CHAN_T(c2s_w_chan_t,logic[AXI_DATA_IN_WIDTH-1:0],logic[AXI_DATA_IN_WIDTH/8-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_B_CHAN_T(c2s_b_chan_t,logic[AXI_ID_IN_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_AR_CHAN_T(c2s_ar_chan_t,logic[AXI_ADDR_WIDTH-1:0],logic[AXI_ID_IN_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_R_CHAN_T(c2s_r_chan_t,logic[AXI_DATA_IN_WIDTH-1:0],logic[AXI_ID_IN_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])

   `AXI_TYPEDEF_REQ_T(c2s_req_t,c2s_aw_chan_t,c2s_w_chan_t,c2s_ar_chan_t)
   `AXI_TYPEDEF_RESP_T(c2s_resp_t,c2s_b_chan_t,c2s_r_chan_t)

   c2s_req_t   dst_req ;
   c2s_resp_t  dst_resp;

   `AXI_TYPEDEF_AW_CHAN_T(s2c_aw_chan_t,logic[AXI_ADDR_WIDTH-1:0],logic[AXI_ID_OUT_S2C_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_W_CHAN_T(s2c_w_chan_t,logic[AXI_DATA_OUT_S2C_WIDTH-1:0],logic[AXI_DATA_OUT_S2C_WIDTH/8-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_B_CHAN_T(s2c_b_chan_t,logic[AXI_ID_OUT_S2C_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_AR_CHAN_T(s2c_ar_chan_t,logic[AXI_ADDR_WIDTH-1:0],logic[AXI_ID_OUT_S2C_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])
   `AXI_TYPEDEF_R_CHAN_T(s2c_r_chan_t,logic[AXI_DATA_OUT_S2C_WIDTH-1:0],logic[AXI_ID_OUT_S2C_WIDTH-1:0],logic[AXI_USER_WIDTH-1:0])

   `AXI_TYPEDEF_REQ_T(s2c_req_t,s2c_aw_chan_t,s2c_w_chan_t,s2c_ar_chan_t)
   `AXI_TYPEDEF_RESP_T(s2c_resp_t,s2c_b_chan_t,s2c_r_chan_t)

   s2c_req_t   src_req ;
   s2c_resp_t  src_resp;

   `AXI_ASSIGN_TO_REQ(src_req,s_data_out_bus)
   `AXI_ASSIGN_FROM_RESP(s_data_out_bus,src_resp)

   // Kill or leave cdc to/from cluster
   if (USE_CLUSTER) begin

     logic s_cluster_isolate_dc;
     logic s_rstn_cluster_sync_soc;

     assign s_rstn_cluster_sync_soc = cluster_rst_ni;

     assign cluster_test_en_o = dft_test_mode_i;
     // isolate dc if the cluster is down
     assign s_cluster_isolate_dc = 1'b0;

     `AXI_ASSIGN_FROM_REQ(s_data_in_bus,dst_req)
     `AXI_ASSIGN_TO_RESP(dst_resp,s_data_in_bus)

     // CLUSTER TO SOC AXI
     axi_cdc_dst #(
       .aw_chan_t (c2s_aw_chan_t),
       .w_chan_t  (c2s_w_chan_t ),
       .b_chan_t  (c2s_b_chan_t ),
       .r_chan_t  (c2s_r_chan_t ),
       .ar_chan_t (c2s_ar_chan_t),
       .axi_req_t (c2s_req_t    ),
       .axi_resp_t(c2s_resp_t   ),
       .LogDepth        ( 3                      )
      ) axi_slave_cdc_i (
       .dst_rst_ni                       ( cluster_rst_ni             ),
       .dst_clk_i                        ( s_soc_clk                  ),
       .dst_req_o                        ( dst_req                    ),
       .dst_resp_i                       ( dst_resp                   ),
       .async_data_slave_aw_wptr_i       ( async_data_slave_aw_wptr_i ),
       .async_data_slave_aw_rptr_o       ( async_data_slave_aw_rptr_o ),
       .async_data_slave_aw_data_i       ( async_data_slave_aw_data_i ),
       .async_data_slave_w_wptr_i        ( async_data_slave_w_wptr_i  ),
       .async_data_slave_w_rptr_o        ( async_data_slave_w_rptr_o  ),
       .async_data_slave_w_data_i        ( async_data_slave_w_data_i  ),
       .async_data_slave_ar_wptr_i       ( async_data_slave_ar_wptr_i ),
       .async_data_slave_ar_rptr_o       ( async_data_slave_ar_rptr_o ),
       .async_data_slave_ar_data_i       ( async_data_slave_ar_data_i ),
       .async_data_slave_b_wptr_o        ( async_data_slave_b_wptr_o  ),
       .async_data_slave_b_rptr_i        ( async_data_slave_b_rptr_i  ),
       .async_data_slave_b_data_o        ( async_data_slave_b_data_o  ),
       .async_data_slave_r_wptr_o        ( async_data_slave_r_wptr_o  ),
       .async_data_slave_r_rptr_i        ( async_data_slave_r_rptr_i  ),
       .async_data_slave_r_data_o        ( async_data_slave_r_data_o  )
      );


    // SOC TO CLUSTER
     axi_cdc_src #(
       .aw_chan_t (s2c_aw_chan_t),
       .w_chan_t  (s2c_w_chan_t),
       .b_chan_t  (s2c_b_chan_t),
       .r_chan_t  (s2c_r_chan_t),
       .ar_chan_t (s2c_ar_chan_t),
       .axi_req_t (s2c_req_t              ),
       .axi_resp_t(s2c_resp_t             ),
      .LogDepth        ( LOG_DEPTH               )
      ) axi_master_cdc_i (
       .src_rst_ni                       ( s_rstn_cluster_sync_soc     ),
       .src_clk_i                        ( s_soc_clk                   ),
       .src_req_i                        ( src_req                     ),
       .src_resp_o                       ( src_resp                    ),
       .async_data_master_aw_wptr_o      ( async_data_master_aw_wptr_o ),
       .async_data_master_aw_rptr_i      ( async_data_master_aw_rptr_i ),
       .async_data_master_aw_data_o      ( async_data_master_aw_data_o ),
       .async_data_master_w_wptr_o       ( async_data_master_w_wptr_o  ),
       .async_data_master_w_rptr_i       ( async_data_master_w_rptr_i  ),
       .async_data_master_w_data_o       ( async_data_master_w_data_o  ),
       .async_data_master_ar_wptr_o      ( async_data_master_ar_wptr_o ),
       .async_data_master_ar_rptr_i      ( async_data_master_ar_rptr_i ),
       .async_data_master_ar_data_o      ( async_data_master_ar_data_o ),
       .async_data_master_b_wptr_i       ( async_data_master_b_wptr_i  ),
       .async_data_master_b_rptr_o       ( async_data_master_b_rptr_o  ),
       .async_data_master_b_data_i       ( async_data_master_b_data_i  ),
       .async_data_master_r_wptr_i       ( async_data_master_r_wptr_i  ),
       .async_data_master_r_rptr_o       ( async_data_master_r_rptr_o  ),
       .async_data_master_r_data_i       ( async_data_master_r_data_i  )
      );

    dc_token_ring_fifo_din #(
        .DATA_WIDTH   ( EVNT_WIDTH   ),
        .BUFFER_DEPTH ( BUFFER_WIDTH )
    ) u_event_dc (
        .clk          ( s_soc_clk               ),
        .rstn         ( s_rstn_cluster_sync_soc ),
        .data         ( s_cl_event_data         ),
        .valid        ( s_cl_event_valid        ),
        .ready        ( s_cl_event_ready        ),
        .write_token  ( cluster_events_wt_o     ),
        .read_pointer ( cluster_events_rp_i     ),
        .data_async   ( cluster_events_da_o     )
    );


    edge_propagator_rx ep_dma_pe_evt_i (
        .clk_i   ( s_soc_clk               ),
        .rstn_i  ( s_rstn_cluster_sync_soc ),
        .valid_o ( s_dma_pe_evt            ),
        .ack_o   ( dma_pe_evt_ack_o        ),
        .valid_i ( dma_pe_evt_valid_i      )
    );

    edge_propagator_rx ep_dma_pe_irq_i (
        .clk_i   ( s_soc_clk               ),
        .rstn_i  ( s_rstn_cluster_sync_soc ),
        .valid_o ( s_dma_pe_irq            ),
        .ack_o   ( dma_pe_irq_ack_o        ),
        .valid_i ( dma_pe_irq_valid_i      )
    );
`ifndef PULP_FPGA_EMUL
    edge_propagator_rx ep_pf_evt_i (
        .clk_i   ( s_soc_clk               ),
        .rstn_i  ( s_rstn_cluster_sync_soc ),
        .valid_o ( s_pf_evt                ),
        .ack_o   ( pf_evt_ack_o            ),
        .valid_i ( pf_evt_valid_i          )
    );
`endif

   end else begin // if (USE_CLUSTER)

     // The AXI slave in the cluster->soc direction is **not** unplugged from the interconnect,
     // because it would require changing the ID width of the exposed AXI port of ControlPULP.
     // Instead, when the cluster is off we tie off this input bus as well.
     assign s_data_in_bus.aw_id = '0;
     assign s_data_in_bus.aw_addr = '0;
     assign s_data_in_bus.aw_len = '0;
     assign s_data_in_bus.aw_size = '0;
     assign s_data_in_bus.aw_burst = '0;
     assign s_data_in_bus.aw_lock = '0;
     assign s_data_in_bus.aw_cache = '0;
     assign s_data_in_bus.aw_prot = '0;
     assign s_data_in_bus.aw_qos = '0;
     assign s_data_in_bus.aw_region = '0;
     assign s_data_in_bus.aw_atop = '0;
     assign s_data_in_bus.aw_user = '0;
     assign s_data_in_bus.aw_valid = '0;
     assign s_data_in_bus.w_data = '0;
     assign s_data_in_bus.w_strb = '0;
     assign s_data_in_bus.w_last = '0;
     assign s_data_in_bus.w_user = '0;
     assign s_data_in_bus.w_valid = '0;
     assign s_data_in_bus.b_ready = '0;
     assign s_data_in_bus.ar_id = '0;
     assign s_data_in_bus.ar_addr = '0;
     assign s_data_in_bus.ar_len = '0;
     assign s_data_in_bus.ar_size = '0;
     assign s_data_in_bus.ar_burst = '0;
     assign s_data_in_bus.ar_lock = '0;
     assign s_data_in_bus.ar_cache = '0;
     assign s_data_in_bus.ar_prot = '0;
     assign s_data_in_bus.ar_qos = '0;
     assign s_data_in_bus.ar_region = '0;
     assign s_data_in_bus.ar_user = '0;
     assign s_data_in_bus.ar_valid = '0;
     assign s_data_in_bus.r_ready = '0;

     assign cluster_events_wt_o = '0;
     assign cluster_events_da_o = '0;

     assign async_data_slave_aw_rptr_o = '0;
     assign async_data_slave_w_rptr_o = '0;
     assign async_data_slave_ar_rptr_o = '0;
     assign async_data_slave_b_wptr_o = '0;
     assign async_data_slave_b_data_o = '0;
     assign async_data_slave_r_wptr_o = '0;
     assign async_data_slave_r_data_o = '0;

     assign async_data_master_aw_wptr_o = '0;
     assign async_data_master_aw_data_o = '0;
     assign async_data_master_ar_wptr_o = '0;
     assign async_data_master_ar_data_o = '0;
     assign async_data_master_w_wptr_o = '0;
     assign async_data_master_w_data_o = '0;
     assign async_data_master_r_rptr_o = '0;
     assign async_data_master_b_rptr_o = '0;

     assign pf_evt_ack_o = '0;
     assign dma_pe_evt_ack_o = '0;
     assign s_dma_pe_evt = '0;
     assign s_dma_pe_irq = '0;
     assign s_pf_evt = '0;
     assign s_cl_event_ready = '0;

     assign cluster_test_en_o = dft_test_mode_i;

     // The AXI master in the soc->cluster direction is terminated with AXI error
     axi_err_slv #(
       .AxiIdWidth  ( AXI_ID_OUT_S2C_WIDTH   ),
       .axi_req_t   ( s2c_req_t              ),
       .axi_resp_t  ( s2c_resp_t             ),
       .Resp        ( axi_pkg::RESP_DECERR   ),
       .ATOPs       ( 1'b0                   ),
       .MaxTrans    ( 4                      )   // Transactions terminate at this slave, so minimize
                                                 // resource consumption by accepting only a few
                                                 // transactions at a time.
     ) i_axi_err_slv (
       .clk_i (s_soc_clk),
       .rst_ni (s_soc_rstn),
       .test_i (1'b0),
       // slave port
       .slv_req_i  ( src_req  ),
       .slv_resp_o ( src_resp )
     );

   end // else: !if(USE_CLUSTER)


    //********************************************************
    //********************* SOC L2 RAM ***********************
    //********************************************************

    // NOTE: The L2 memories are outside the control-pulp module!

    //********************************************************
    //******              SOC BOOT ROM             ***********
    //********************************************************

    boot_rom #(
        .ROM_ADDR_WIDTH(ROM_ADDR_WIDTH),
        .MACRO_ROM(MACRO_ROM)
    ) boot_rom_i (
        .clk_i       ( s_soc_clk       ),
        .rst_ni      ( s_soc_rstn      ),
        .init_ni     ( 1'b1            ),
        .mem_slave   ( s_mem_rom_bus   ),
        .test_mode_i ( dft_test_mode_i )
    );

    //********************************************************
    //********************* SOC PERIPHERALS ******************
    //********************************************************

    soc_peripherals #(
        .CORE_TYPE          ( CORE_TYPE                             ),
        .MEM_ADDR_WIDTH     ( L2_MEM_ADDR_WIDTH+$clog2(N_L2_BANKS)  ),
        .APB_ADDR_WIDTH     ( 32                                    ),
        .APB_DATA_WIDTH     ( 32                                    ),
        .NB_CORES           ( NB_CORES                              ),
        .NB_CLUSTERS        ( `NB_CLUSTERS                          ),
        .EVNT_WIDTH         ( EVNT_WIDTH                            ),
        .NGPIO              ( NGPIO                                 ),
        .NBIT_PADCFG        ( NBIT_PADCFG                           ),
        .N_UART             ( N_UART                                ),
        .N_SPI              ( N_SPI                                 ),
        .N_I2C              ( N_I2C                                 ),
        .N_I2C_SLV          ( N_I2C_SLV                             ),
        .SIM_STDOUT         ( SIM_STDOUT                            ),

        // AXI widths for spi_slv, i2c_slvs AXI conversion within soc_peripherals
        .AXI_ADDR_WIDTH     ( AXI_ADDR_WIDTH                        ),
        .AXI_DATA_IN_WIDTH  ( 32                                    ),
        .AXI_ID_IN_WIDTH    ( AXI_ID_IN_WIDTH                       ),
        .AXI_USER_WIDTH     ( AXI_USER_WIDTH                        )

    ) soc_peripherals_i (

        .clk_i                  ( s_soc_clk              ),
        .periph_clk_i,
        .rst_ni                 ( s_soc_rstn             ),
        .sel_clk_i              ( s_sel_clk              ),
        .slow_clk_i             ( ref_clk_i              ),

        .dft_test_mode_i,
        .dft_cg_enable_i,

        .bootsel_valid_i        ( bootsel_valid_i        ),
        .bootsel_i              ( bootsel_i              ),

        .fc_fetch_en_valid_i    ( fc_fetch_en_valid_i    ),
        .fc_fetch_en_i          ( fc_fetch_en_i          ),

        .fc_bootaddr_o          ( s_fc_bootaddr          ),
        .fc_fetchen_o           ( s_fc_fetchen           ),

        .apb_slave              ( s_apb_periph_bus       ),

        .apb_eu_master          ( s_apb_eu_bus           ),
        .apb_clic_master        ( s_apb_clic_bus         ),
        .apb_debug_master       ( s_apb_debug_bus        ),
        .apb_hwpe_master        ( s_apb_hwpe_bus         ),
        .apb_serial_link_master ( apb_serial_link_bus    ),
        .apb_clk_ctrl_master    ( apb_clk_ctrl_bus       ),
        .apb_pad_cfg_master     ( apb_pad_cfg_bus        ),
        .apb_sdma_cfg_master    ( s_apb_sdma_bus         ),

        .l2_rx_master           ( s_lint_udma_rx_bus     ),
        .l2_tx_master           ( s_lint_udma_tx_bus     ),

        .axi_mst_spi_slv        ( s_axi_spi              ),

        .soc_jtag_reg_i         ( soc_jtag_reg_tap       ),
        .soc_jtag_reg_o         ( soc_jtag_reg_soc       ),

        .fc_hwpe_events_i       ( s_fc_hwpe_events       ),
        .fc_events_o            ( s_fc_events            ),

        .dma_pe_evt_i           ( s_dma_pe_evt           ),
        .dma_pe_irq_i           ( s_dma_pe_irq           ),
        .pf_evt_i               ( s_pf_evt               ),

        .gpio_in                ( gpio_in_i              ),
        .gpio_out               ( gpio_out_o             ),
        .gpio_dir               ( gpio_dir_o             ),
        .gpio_padcfg            ( gpio_cfg_o             ),

        //UART
        .uart_tx                ( uart_tx_o              ),
        .uart_rx                ( uart_rx_i              ),

        //I2C
        .i2c_scl_i              ( i2c_scl_i              ),
        .i2c_scl_o              ( i2c_scl_o              ),
        .i2c_scl_oe_o           ( i2c_scl_oe_o           ),
        .i2c_sda_i              ( i2c_sda_i              ),
        .i2c_sda_o              ( i2c_sda_o              ),
        .i2c_sda_oe_o           ( i2c_sda_oe_o           ),

        //I2C slave
        .i2c_slv_scl_i          ( i2c_slv_scl_i          ),
        .i2c_slv_scl_o          ( i2c_slv_scl_o          ),
        .i2c_slv_scl_oe_o       ( i2c_slv_scl_oe_o       ),
        .i2c_slv_sda_i          ( i2c_slv_sda_i          ),
        .i2c_slv_sda_o          ( i2c_slv_sda_o          ),
        .i2c_slv_sda_oe_o       ( i2c_slv_sda_oe_o       ),

         //SPI MASTER
        .spi_clk_o              ( spi_clk_o              ),
        .spi_csn_o              ( spi_csn_o              ),
        .spi_oen_o              ( spi_oen_o              ),
        .spi_sdo_o              ( spi_sdo_o              ),
        .spi_sdi_i              ( spi_sdi_i              ),

         //SPI SLAVE
        .spi_clk_i              ( spi_clk_i              ),
        .spi_csn_i              ( spi_csn_i              ),
        .spi_oen_slv_o          ( spi_oen_slv_o          ),
        .spi_sdo_slv_o          ( spi_sdo_slv_o          ),
        .spi_sdi_slv_i          ( spi_sdi_slv_i          ),

        //INTER-SOCKET MUX SIGNALS
        .sel_spi_dir_o          ( sel_spi_dir_o          ),
        .sel_i2c_mux_o          ( sel_i2c_mux_o          ),

        .timer_ch0_o            ( timer_ch0_o            ),
        .timer_ch1_o            ( timer_ch1_o            ),
        .timer_ch2_o            ( timer_ch2_o            ),
        .timer_ch3_o            ( timer_ch3_o            ),

        .cl_event_data_o        ( s_cl_event_data        ),
        .cl_event_valid_o       ( s_cl_event_valid       ),
        .cl_event_ready_i       ( s_cl_event_ready       ),

        .fc_event_data_o        ( s_fc_event_data        ),
        .fc_event_valid_o       ( s_fc_event_valid       ),
        .fc_event_ready_i       ( s_fc_event_ready       ),

        .cluster_pow_o          ( cluster_pow_o          ),
        .cluster_byp_o          ( cluster_byp_o          ),
        .cluster_boot_addr_o    ( cluster_boot_addr_o    ),
        .cluster_fetch_enable_o ( cluster_fetch_enable_o ),
        .cluster_rstn_o         ( cluster_rst_reg_no     ),
        .cluster_irq_o          ( cluster_irq_o          ),

        .wdt_alert_o,
        .wdt_alert_clear_i,

        .bus_instr_err_i        ( s_lint_fc_instr_bus.r_opc & s_lint_fc_instr_bus.r_valid ),
        .bus_data_err_i         ( s_lint_fc_data_bus.r_opc  & s_lint_fc_data_bus.r_valid  ),

        .axi_i2c_slv_bmc        ( axi_i2c_slv_bmc        ),
        .axi_i2c_slv_1          ( axi_i2c_slv_1          )
    );


    fc_subsystem #(
        .CORE_TYPE  ( CORE_TYPE          ),
        .PULP_XPULP ( PULP_XPULP         ),
        .USE_FPU    ( USE_FPU            ),
        .ZFINX      ( ZFINX              ),
        .N_EXT_PERF_COUNTERS( N_PERF_COUNTERS ),
        .CORE_ID    ( FC_CORE_CORE_ID    ),
        .CLUSTER_ID ( FC_CORE_CLUSTER_ID ),
        .USE_HWPE   ( USE_HWPE           ),
        .NUM_INTERRUPTS ( NUM_INTERRUPTS )
    ) fc_subsystem_i (
        .clk_i               ( s_soc_clk                     ),
        .rst_ni              ( s_soc_rstn                    ),

        .test_en_i           ( dft_test_mode_i               ),

        .boot_addr_i         ( s_fc_bootaddr                 ),

        .fetch_en_i          ( s_fc_fetchen                  ),

        .l2_data_master      ( s_lint_fc_data_bus            ),
        .l2_instr_master     ( s_lint_fc_instr_bus           ),
        .l2_shadow_master    ( s_lint_fc_shadow_bus          ),
        .l2_hwpe_master      ( s_lint_hwpe_bus               ),
        .apb_slave_eu        ( s_apb_eu_bus                  ),
        .apb_slave_clic      ( s_apb_clic_bus                ),
        .apb_slave_hwpe      ( s_apb_hwpe_bus                ),
        .debug_req_i         ( dm_debug_req[FC_CORE_MHARTID] ),

        .event_fifo_valid_i  ( s_fc_event_valid              ),
        .event_fifo_fulln_o  ( s_fc_event_ready              ),
        .event_fifo_data_i   ( s_fc_event_data               ),
        .events_i            ( s_fc_events                   ),

        .hwpe_events_o       ( s_fc_hwpe_events              ),

        // SDMA events
        .sdma_term_event_i   ( s_sdma_term_event             ),
        .sdma_busy_i         ( s_sdma_busy                   ),

        .supervisor_mode_o   ( s_supervisor_mode             ),

        // External interrupts
        .scg_irq_i,
        .scp_irq_i,
        .scp_secure_irq_i,
        .mbox_irq_i,
        .mbox_secure_irq_i
    );

    // Sensor DMA

    // Configuration parameters
    localparam int unsigned SDMA_NB_OUTSND_BURSTS = 8;
    localparam int unsigned SDMA_REG_DATA_WIDTH = 32;
    localparam int unsigned SDMA_REG_ADDR_WIDTH = 32;

    dmac_wrap_fc_idma #(
      .AXI_ADDR_WIDTH   ( AXI_ADDR_WIDTH      ),
      .AXI_DATA_WIDTH   ( AXI_DATA_OUT_S2E_WIDTH ),
      .AXI_USER_WIDTH   ( AXI_USER_WIDTH      ),
      .AXI_ID_WIDTH_MST_1 ( AXI_ID_OUT_S2C_WIDTH), // to ext ID
      .AXI_ID_WIDTH_MST_2 ( AXI_ID_IN_WIDTH   ), // to tcdm ID
      .DATA_WIDTH       ( SDMA_REG_DATA_WIDTH ),
      .ADDR_WIDTH       ( SDMA_REG_ADDR_WIDTH ),
      .NUM_STREAMS      ( 1                   ),
      .L2_SIZE          ( L2_SIZE             ), // size of src/dst memory
      .NB_OUTSND_BURSTS ( SDMA_NB_OUTSND_BURSTS )
    ) i_sensor_dma (
      .clk_i           (s_soc_clk                       ),
      .rst_ni          (s_soc_rstn                      ),
      .test_mode_i     (dft_test_mode_i                 ),
      .apb_sdma_cfg_bus(s_apb_sdma_bus),
      .axi_tcdm_master (s_axi_tcdm_sdma_mst),
      .axi_ext_master  (s_axi_ext_sdma_mst),
      .term_event_o    (s_sdma_term_event), // to clic
      .term_irq_o      (), // unused for now
      .busy_o          (s_sdma_busy)  // to clic
    );

    // Upsize AXI data width SOC->EXT (32b->64b) direction in the core path
    // This is needed for compliance with the 64b DMA coupled with the core, that
    // can handle 64b transfers without the mem->axi bottleneck (DW = 32b) of the core
    // The two 64b ports (1 from the core, 1 from the sdma) are muxed to the unique 64b output port

    axi_dw_converter_intf #(
      .AXI_ID_WIDTH            ( AXI_ID_OUT_S2C_WIDTH),
      .AXI_ADDR_WIDTH          ( AXI_ADDR_WIDTH     ),
      .AXI_SLV_PORT_DATA_WIDTH ( AXI_DATA_OUT_S2C_WIDTH ), //32b
      .AXI_MST_PORT_DATA_WIDTH ( AXI_DATA_OUT_S2E_WIDTH ), //64b
      .AXI_USER_WIDTH          ( AXI_USER_WIDTH     ),
      .AXI_MAX_READS           ( 1                  )
    ) axi_dw_upsize_32_64_i (
      .clk_i  ( s_soc_clk       ),
      .rst_ni ( s_soc_rstn      ),
      .slv    ( s_axi_ext_core_mst ),
      .mst    ( s_axi_ext_core_dw_mst )
    );
    
    // Arbitrate between core and sdma to communicate with the single external port
    axi_mux_intf #(
      .SLV_AXI_ID_WIDTH( AXI_ID_OUT_S2C_WIDTH ),
      .MST_AXI_ID_WIDTH( AXI_ID_OUT_S2E_WIDTH ),
      .AXI_ADDR_WIDTH( AXI_ADDR_WIDTH     ),
      .AXI_DATA_WIDTH( AXI_DATA_OUT_S2E_WIDTH ),
      .AXI_USER_WIDTH( AXI_USER_WIDTH     ),
      .NO_SLV_PORTS( 2 ),
      .MAX_W_TRANS( 1 ),
      .FALL_THROUGH( 1'b1 )
    ) i_axi64_ext_mux (
      .clk_i(s_soc_clk),
      .rst_ni(s_soc_rstn),
      .test_i(dft_test_mode_i),
      .slv(axi_mux_ext_slv),
      .mst(axi_ext_mst)
    );

    // FC interconnect
    soc_interconnect_wrap #(
        .NR_HWPE_PORTS       ( NB_HWPE_PORTS    ),
        .NR_L2_PORTS         ( N_L2_BANKS       ),
        .AXI_USER_WIDTH      ( AXI_USER_WIDTH   ),
        .AXI_IN_ID_WIDTH     ( AXI_ID_IN_WIDTH  ),
        .N_EXT_MASTERS_TO_SOC( N_EXT_MASTERS_TO_SOC ),
        .N_EXT_MASTERS_TO_SOC_PERIPH( N_EXT_MASTERS_TO_SOC_PERIPH)
    ) i_soc_interconnect_wrap (
        .clk_i            ( s_soc_clk            ),
        .rst_ni           ( s_soc_rstn           ),
        .test_en_i        ( dft_test_mode_i      ),
        .tcdm_fc_data     ( s_lint_fc_data_bus   ),
        .tcdm_fc_instr    ( s_lint_fc_instr_bus  ),
        .tcdm_fc_shadow   ( s_lint_fc_shadow_bus ),
        .tcdm_udma_rx     ( s_lint_udma_rx_bus   ),
        .tcdm_udma_tx     ( s_lint_udma_tx_bus   ),
        .tcdm_debug       ( s_lint_debug_bus     ),
        .tcdm_hwpe        ( s_lint_hwpe_bus      ),

        // ext-to-pms direction (wrapped interface)
        .axi_master_plug  ( ext_masters_to_soc  ), // from external in-band modules (cluster, ext)
        .axi_master_plug_periph  ( ext_masters_to_soc_periph  ), // from external out-of-band periph (spi, i2c_1, i2c_2)

        // pms-to-ext direction (discrete interfaces)
        .axi_slave_plug   ( s_data_out_bus      ), // to_cluster
        .axi_ext_mst      ( s_axi_ext_core_mst  ), // to ext
        .apb_peripheral_bus    ( s_apb_periph_bus        ), // to apb_periph

        .l2_interleaved_slaves ( s_mem_l2_bus            ), // to interleaved L2
        .l2_private_slaves     ( s_mem_l2_pri_bus        ), // to private L2
        .boot_rom_slave        ( s_mem_rom_bus           )  // to bootrom
    );

    // Debug Subsystem
    dmi_jtag #(
        .IdcodeValue          ( `DMI_JTAG_IDCODE    )
    ) i_dmi_jtag (
        .clk_i                ( s_soc_clk           ),
        .rst_ni               ( s_soc_rstn          ),
        .testmode_i           ( dft_test_mode_i     ),
        .dmi_req_o            ( jtag_dmi_req        ),
        .dmi_req_valid_o      ( jtag_req_valid      ),
        .dmi_req_ready_i      ( debug_req_ready     ),
        .dmi_resp_i           ( debug_resp          ),
        .dmi_resp_ready_o     ( jtag_resp_ready     ),
        .dmi_resp_valid_i     ( jtag_resp_valid     ),
        .dmi_rst_no           (                     ), // not connected
        .tck_i                ( jtag_tck_i          ),
        .tms_i                ( jtag_tms_i          ),
        .trst_ni              ( jtag_trst_ni        ),
        .td_i                 ( jtag_tdi_i          ),
        .td_o                 ( int_td              ),
        .tdo_oe_o             (                     )
    );

    // set hartinfo
    always_comb begin: set_hartinfo
        for (int hartid = 0; hartid < NrHarts; hartid = hartid + 1) begin
            hartinfo[hartid] = RI5CY_HARTINFO;
        end
    end

    // redirect debug request from dm to correct cluster core
    for (genvar dbg_var = 0; dbg_var < NB_CORES; dbg_var = dbg_var + 1) begin : gen_debug_valid
        assign cluster_dbg_irq_valid_o[dbg_var] = dm_debug_req[cluster_core_id[dbg_var]];
    end

    dm_top #(
       .NrHarts           ( NrHarts                   ),
       .BusWidth          ( 32                        ),
       .ReadByteEnable    ( 0                         ),
       .SelectableHarts   ( SELECTABLE_HARTS          )
    ) i_dm_top (

       .clk_i             ( s_soc_clk                 ),
       .rst_ni            ( s_soc_rstn                ),
       .testmode_i        ( 1'b0                      ),
       .ndmreset_o        (                           ),
       .dmactive_o        (                           ), // active debug session
       .debug_req_o       ( dm_debug_req              ),
       .unavailable_i     ( ~SELECTABLE_HARTS         ),
       .hartinfo_i        ( hartinfo                  ),

       .slave_req_i       ( slave_req                 ),
       .slave_we_i        ( slave_we                  ),
       .slave_addr_i      ( slave_addr                ),
       .slave_be_i        ( slave_be                  ),
       .slave_wdata_i     ( slave_wdata               ),
       .slave_rdata_o     ( slave_rdata               ),

       .master_req_o      ( s_lint_riscv_jtag_bus.req      ),
       .master_add_o      ( s_lint_riscv_jtag_bus.add      ),
       .master_we_o       ( lint_riscv_jtag_bus_master_we  ),
       .master_wdata_o    ( s_lint_riscv_jtag_bus.wdata    ),
       .master_be_o       ( s_lint_riscv_jtag_bus.be       ),
       .master_gnt_i      ( s_lint_riscv_jtag_bus.gnt      ),
       .master_r_valid_i  ( s_lint_riscv_jtag_bus.r_valid  ),
       .master_r_rdata_i  ( s_lint_riscv_jtag_bus.r_rdata  ),
       .master_r_other_err_i ('0                           ),
       .master_r_err_i       ('0                           ),

       .dmi_rst_ni        ( s_soc_rstn                ),
       .dmi_req_valid_i   ( jtag_req_valid            ),
       .dmi_req_ready_o   ( debug_req_ready           ),
       .dmi_req_i         ( jtag_dmi_req              ),
       .dmi_resp_valid_o  ( jtag_resp_valid           ),
       .dmi_resp_ready_i  ( jtag_resp_ready           ),
       .dmi_resp_o        ( debug_resp                )
    );
    assign s_lint_riscv_jtag_bus.wen = ~lint_riscv_jtag_bus_master_we;

    jtag_tap_top  #(
        .IDCODE_VALUE             ( `PULP_JTAG_IDCODE   )
    ) jtag_tap_top_i (
        .tck_i                    ( jtag_tck_i         ),
        .trst_ni                  ( jtag_trst_ni       ),
        .tms_i                    ( jtag_tms_i         ),
        .td_i                     ( int_td             ),
        .td_o                     ( jtag_tdo_o         ),

        .test_clk_i               ( 1'b0               ),
        .test_rstn_i              ( s_soc_rstn         ),

        .jtag_shift_dr_o          ( s_jtag_shift_dr    ),
        .jtag_update_dr_o         ( s_jtag_update_dr   ),
        .jtag_capture_dr_o        ( s_jtag_capture_dr  ),

        .axireg_sel_o             ( s_jtag_axireg_sel  ),
        .dbg_axi_scan_in_o        ( s_jtag_axireg_tdi  ),
        .dbg_axi_scan_out_i       ( s_jtag_axireg_tdo  ),
        .soc_jtag_reg_i           ( soc_jtag_reg_soc   ),
        .soc_jtag_reg_o           ( soc_jtag_reg_tap   ),
        .sel_clk_o                ( s_sel_clk          )
    );

    lint_jtag_wrap i_lint_jtag (
        .tck_i                    ( jtag_tck_i           ),
        .tdi_i                    ( s_jtag_axireg_tdi    ),
        .trstn_i                  ( jtag_trst_ni         ),
        .tdo_o                    ( s_jtag_axireg_tdo    ),
        .shift_dr_i               ( s_jtag_shift_dr      ),
        .pause_dr_i               ( 1'b0                 ),
        .update_dr_i              ( s_jtag_update_dr     ),
        .capture_dr_i             ( s_jtag_capture_dr    ),
        .lint_select_i            ( s_jtag_axireg_sel    ),
        .clk_i                    ( s_soc_clk            ),
        .rst_ni                   ( s_soc_rstn           ),
        .jtag_lint_master         ( s_lint_pulp_jtag_bus )
    );

    tcdm_arbiter_2x1 jtag_lint_arbiter_i
     (
        .clk_i(s_soc_clk),
        .rst_ni(s_soc_rstn),
        .tcdm_bus_1_i(s_lint_riscv_jtag_bus),
        .tcdm_bus_0_i(s_lint_pulp_jtag_bus),
        .tcdm_bus_o(s_lint_debug_bus)
    );

    apb2per #(
        .PER_ADDR_WIDTH ( 32  ),
        .APB_ADDR_WIDTH ( 32  )
    ) apb2per_newdebug_i (
        .clk_i                ( s_soc_clk               ),
        .rst_ni               ( s_soc_rstn              ),

        .PADDR                ( s_apb_debug_bus.paddr   ),
        .PWDATA               ( s_apb_debug_bus.pwdata  ),
        .PWRITE               ( s_apb_debug_bus.pwrite  ),
        .PSEL                 ( s_apb_debug_bus.psel    ),
        .PENABLE              ( s_apb_debug_bus.penable ),
        .PRDATA               ( s_apb_debug_bus.prdata  ),
        .PREADY               ( s_apb_debug_bus.pready  ),
        .PSLVERR              ( s_apb_debug_bus.pslverr ),

        .per_master_req_o     ( slave_req               ),
        .per_master_add_o     ( slave_addr              ),
        .per_master_we_o      ( slave_we                ),
        .per_master_wdata_o   ( slave_wdata             ),
        .per_master_be_o      ( slave_be                ),
        .per_master_gnt_i     ( slave_grant             ),
        .per_master_r_valid_i ( slave_valid             ),
        .per_master_r_opc_i   ( '0                      ),
        .per_master_r_rdata_i ( slave_rdata             )
     );

     assign slave_grant = slave_req;
     always_ff @(posedge s_soc_clk or negedge s_soc_rstn) begin : apb2per_valid
         if(~s_soc_rstn) begin
             slave_valid <= 0;
         end else begin
             slave_valid <= slave_grant;
         end
     end

endmodule

// Local Variables:
// verilog-indent-level: 4
// verilog-indent-level-module: 4
// verilog-indent-level-declaration: 4
// verilog-indent-level-behavioral: 4
// verilog-case-indent: 4
// verilog-cexp-indent: 4
// End:
